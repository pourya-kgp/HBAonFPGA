----------------------------------------------------------------------------------------------------
-- Author           : Pourya Khodagholipour (P.KH)
-- Project Name     : HBA (Hardware Bee Algorithm)
-- File Name        : TSP_Dist_One_Port_ROM_Sync
-- Module Name      : TSP_Dist_One_Port_ROM_Sync
-- HDL Standard     : VHDL
-- Approach         : Behavioral
-- Description      : Single-port ROM with synchronous read (Block RAM)
-- Comments         : berlin52 Database Distance matrix
-- Dependencies     : ---
-- Target Devices   : Virtex 5 - XC5VLX330
-- Speed Estimation : ---
-- Area  Estimation : 2 RAM/FIFO
-- Tools            : ISE Design Suite v14.7 - Altera Quartus 16.1 Lite
-- Module Version   : 
-- Creation Date    : 2016/08
-- Revision Date    : 2024/07/08
----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity TSP_Dist_One_Port_ROM_Sync is
	generic (
				ADDR_WIDTH : natural := 11;
				DATA_WIDTH : natural := 32);
	port    (
				CLK        : in  std_logic;
				ADDR       : in  std_logic_vector (ADDR_WIDTH-1 downto 0);
				DATA       : out std_logic_vector (DATA_WIDTH-1 downto 0));
end TSP_Dist_One_Port_ROM_Sync;

architecture Behavioral of TSP_Dist_One_Port_ROM_Sync is

	type ROM_Type is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector (DATA_WIDTH-1 downto 0);
	constant ROM : ROM_Type := (
			"11111111111111111111111111111111" , -- ADDR 0
			"00000000000010100010100111111100" , -- ADDR 1
			"00000000000001000100101000011010" , -- ADDR 2
			"00000000000001100000100101010001" , -- ADDR 3
			"00000000000001000111000110000100" , -- ADDR 4
			"00000000000001001111101001111011" , -- ADDR 5
			"00000000000010011100011100100000" , -- ADDR 6
			"00000000000001101000001101111110" , -- ADDR 7
			"00000000000010010010100001111011" , -- ADDR 8
			"00000000000010001001000100111111" , -- ADDR 9
			"00000000000011111110001001001101" , -- ADDR 10
			"00000000000010011111111010101011" , -- ADDR 11
			"00000000000011101110000010011000" , -- ADDR 12
			"00000000000100010001101000000010" , -- ADDR 13
			"00000000000001001001000000100000" , -- ADDR 14
			"00000000000000111111011111010000" , -- ADDR 15
			"00000000000001101000110111011111" , -- ADDR 16
			"00000000000000100111011100010011" , -- ADDR 17
			"00000000000001001010011101101000" , -- ADDR 18
			"00000000000000110011010010001100" , -- ADDR 19
			"00000000000001000110000011001011" , -- ADDR 20
			"00000000000000001011010000010010" , -- ADDR 21
			"00000000000000101100001110111001" , -- ADDR 22
			"00000000000001000011000010011111" , -- ADDR 23
			"00000000000001100100000110101110" , -- ADDR 24
			"00000000000010110001111110001100" , -- ADDR 25
			"00000000000011000010111100110010" , -- ADDR 26
			"00000000000010101100100110111001" , -- ADDR 27
			"00000000000001100011001011110111" , -- ADDR 28
			"00000000000001010111111010000101" , -- ADDR 29
			"00000000000000100011101111000101" , -- ADDR 30
			"00000000000000010110000110111010" , -- ADDR 31
			"00000000000011001001111110110011" , -- ADDR 32
			"00000000000000100000111110110101" , -- ADDR 33
			"00000000000000011101101100110111" , -- ADDR 34
			"00000000000000011110100001001000" , -- ADDR 35
			"00000000000000110010110001011110" , -- ADDR 36
			"00000000000000111010101100100000" , -- ADDR 37
			"00000000000000101000100101000000" , -- ADDR 38
			"00000000000000110011000000011110" , -- ADDR 39
			"00000000000001100000100001110100" , -- ADDR 40
			"00000000000010001010001000100100" , -- ADDR 41
			"00000000000001110001001111001000" , -- ADDR 42
			"00000000000000100101101101000010" , -- ADDR 43
			"00000000000000111010101001010000" , -- ADDR 44
			"00000000000001000100010100111010" , -- ADDR 45
			"00000000000011000001001011110001" , -- ADDR 46
			"00000000000001000001010000100101" , -- ADDR 47
			"00000000000000001111101000011111" , -- ADDR 48
			"00000000000000110100111111111011" , -- ADDR 49
			"00000000000011000000101110000111" , -- ADDR 50
			"00000000000100101001111101101101" , -- ADDR 51
			"00000000000010011110100001101111" , -- ADDR 52
			"00000000000011111111101000110011" , -- ADDR 53
			"00000000000011100110101111111001" , -- ADDR 54
			"00000000000011101110110010100101" , -- ADDR 55
			"00000000000000001010111111001000" , -- ADDR 56
			"00000000000011101001011011110111" , -- ADDR 57
			"00000000000100010101000101101100" , -- ADDR 58
			"00000000000100010100100110110111" , -- ADDR 59
			"00000000000110010000000110000100" , -- ADDR 60
			"00000000000100110011010001011110" , -- ADDR 61
			"00000000000101011111100101001110" , -- ADDR 62
			"00000000000101110010000011001110" , -- ADDR 63
			"00000000000011101001110101111111" , -- ADDR 64
			"00000000000010110000110001000010" , -- ADDR 65
			"00000000000001111000110010110101" , -- ADDR 66
			"00000000000010010001011000011011" , -- ADDR 67
			"00000000000011001101111010001001" , -- ADDR 68
			"00000000000010001001110011110101" , -- ADDR 69
			"00000000000001011111110100001100" , -- ADDR 70
			"00000000000010011011011000000000" , -- ADDR 71
			"00000000000001111100011110000100" , -- ADDR 72
			"00000000000011100001000011000000" , -- ADDR 73
			"00000000000011111011001011101110" , -- ADDR 74
			"00000000000100100010111001011000" , -- ADDR 75
			"00000000000100111101110000000101" , -- ADDR 76
			"00000000000100101111101001001100" , -- ADDR 77
			"00000000000010011011000010001100" , -- ADDR 78
			"00000000000001011111010100110000" , -- ADDR 79
			"00000000000010000100001000101001" , -- ADDR 80
			"00000000000010110010001110010000" , -- ADDR 81
			"00000000000101101011011101000011" , -- ADDR 82
			"00000000000010111110111100000001" , -- ADDR 83
			"00000000000010111101101100010101" , -- ADDR 84
			"00000000000010111111101001101000" , -- ADDR 85
			"00000000000011010001011001100100" , -- ADDR 86
			"00000000000011011010111110101011" , -- ADDR 87
			"00000000000011001010001000111100" , -- ADDR 88
			"00000000000011010100010101101101" , -- ADDR 89
			"00000000000011011010110010101100" , -- ADDR 90
			"00000000000000011001000010111111" , -- ADDR 91
			"00000000000100010010010101111110" , -- ADDR 92
			"00000000000010110101110110110011" , -- ADDR 93
			"00000000000011001000111111110110" , -- ADDR 94
			"00000000000011010001101111001100" , -- ADDR 95
			"00000000000100011001000100100111" , -- ADDR 96
			"00000000000011011110001111011110" , -- ADDR 97
			"00000000000010110001101111001011" , -- ADDR 98
			"00000000000010010001100100100011" , -- ADDR 99
			"00000000000101011011000011110101" , -- ADDR 100
			"00000000000110100010111101010001" , -- ADDR 101
			"00000000000010010011010101110111" , -- ADDR 102
			"00000000000001111100010000010001" , -- ADDR 103
			"00000000000010000100011100110101" , -- ADDR 104
			"00000000000010010101000100001110" , -- ADDR 105
			"00000000000001001011001101011010" , -- ADDR 106
			"00000000000001110110100100001100" , -- ADDR 107
			"00000000000001110110111101011111" , -- ADDR 108
			"00000000000100110101010000000001" , -- ADDR 109
			"00000000000011011001100111100001" , -- ADDR 110
			"00000000000100110000101000001110" , -- ADDR 111
			"00000000000101010101101110110100" , -- ADDR 112
			"00000000000001111011010000101100" , -- ADDR 113
			"00000000000010000011001100111001" , -- ADDR 114
			"00000000000000110101000011100001" , -- ADDR 115
			"00000000000000100000110111100101" , -- ADDR 116
			"00000000000000110010100010011010" , -- ADDR 117
			"00000000000001101011101010000101" , -- ADDR 118
			"00000000000001000110011100010011" , -- ADDR 119
			"00000000000000111010101110001000" , -- ADDR 120
			"00000000000001011000001011011011" , -- ADDR 121
			"00000000000001111011011101011101" , -- ADDR 122
			"00000000000010011111010011110110" , -- ADDR 123
			"00000000000011110101100101111001" , -- ADDR 124
			"00000000000100000100101001110110" , -- ADDR 125
			"00000000000011101100111001010010" , -- ADDR 126
			"00000000000010011110111111110001" , -- ADDR 127
			"00000000000001111011000110001111" , -- ADDR 128
			"00000000000000110011000000011110" , -- ADDR 129
			"00000000000000111011110111010100" , -- ADDR 130
			"00000000000011011100100011100100" , -- ADDR 131
			"00000000000001100000000110000101" , -- ADDR 132
			"00000000000001011011001110100000" , -- ADDR 133
			"00000000000001011001110001010000" , -- ADDR 134
			"00000000000001101101001111101001" , -- ADDR 135
			"00000000000001110000110100001000" , -- ADDR 136
			"00000000000001011111110000101101" , -- ADDR 137
			"00000000000001101000001101111110" , -- ADDR 138
			"00000000000000111100010011000110" , -- ADDR 139
			"00000000000010000110010011001011" , -- ADDR 140
			"00000000000010000111111000110101" , -- ADDR 141
			"00000000000001101010000000010011" , -- ADDR 142
			"00000000000000110101101010110101" , -- ADDR 143
			"00000000000010000110111011100011" , -- ADDR 144
			"00000000000100000101110010110111" , -- ADDR 145
			"00000000000001111011001111100010" , -- ADDR 146
			"00000000000001000110011011100111" , -- ADDR 147
			"00000000000001110001000110010001" , -- ADDR 148
			"00000000000011110010111111110010" , -- ADDR 149
			"00000000000101101010001101001010" , -- ADDR 150
			"00000000000000011001011111010011" , -- ADDR 151
			"00000000000000010001000000001010" , -- ADDR 152
			"00000000000011111010100100111101" , -- ADDR 153
			"00000000000010000000001011001000" , -- ADDR 154
			"00000000000010010101001010111011" , -- ADDR 155
			"00000000000010000010010110001101" , -- ADDR 156
			"00000000000010100001111010011001" , -- ADDR 157
			"00000000000001000111110111011100" , -- ADDR 158
			"00000000000010101101100110100001" , -- ADDR 159
			"00000000000011011010111111110001" , -- ADDR 160
			"00000000000000011000011100011101" , -- ADDR 161
			"00000000000001011101110011011100" , -- ADDR 162
			"00000000000011000011010111111010" , -- ADDR 163
			"00000000000010000001111110000001" , -- ADDR 164
			"00000000000001110011111000111100" , -- ADDR 165
			"00000000000001111010001110010001" , -- ADDR 166
			"00000000000010100110011000001111" , -- ADDR 167
			"00000000000001101010100101111110" , -- ADDR 168
			"00000000000010000011010001100111" , -- ADDR 169
			"00000000000000011110100101110100" , -- ADDR 170
			"00000000000000011010101010010010" , -- ADDR 171
			"00000000000001111110000010001100" , -- ADDR 172
			"00000000000010000000100111010110" , -- ADDR 173
			"00000000000001100101111010011001" , -- ADDR 174
			"00000000000010001101100100011111" , -- ADDR 175
			"00000000000010101000010101111001" , -- ADDR 176
			"00000000000010000100000010111000" , -- ADDR 177
			"00000000000001011010011101101100" , -- ADDR 178
			"00000000000001111110010011100101" , -- ADDR 179
			"00000000000001000001000100111000" , -- ADDR 180
			"00000000000001000011001011000000" , -- ADDR 181
			"00000000000001000010000100001001" , -- ADDR 182
			"00000000000000101110011110111010" , -- ADDR 183
			"00000000000000100101111001101010" , -- ADDR 184
			"00000000000000111000010001011001" , -- ADDR 185
			"00000000000000101101111101111010" , -- ADDR 186
			"00000000000010000100111100011101" , -- ADDR 187
			"00000000000011101000000000111001" , -- ADDR 188
			"00000000000000111011110111010100" , -- ADDR 189
			"00000000000001001010111100111010" , -- ADDR 190
			"00000000000001100100010111011000" , -- ADDR 191
			"00000000000000111000010100110001" , -- ADDR 192
			"00000000000010100001000001101100" , -- ADDR 193
			"00000000000000100001100001001111" , -- ADDR 194
			"00000000000001010100010010100110" , -- ADDR 195
			"00000000000001110100100110111000" , -- ADDR 196
			"00000000000001100000111011011100" , -- ADDR 197
			"00000000000011011101110101011111" , -- ADDR 198
			"00000000000000001000101000011011" , -- ADDR 199
			"00000000000011100001011111001010" , -- ADDR 200
			"00000000000001110010111000011110" , -- ADDR 201
			"00000000000010001110011111001111" , -- ADDR 202
			"00000000000001111101010110111101" , -- ADDR 203
			"00000000000010111001101111100101" , -- ADDR 204
			"00000000000001011101010111011010" , -- ADDR 205
			"00000000000010111011110000010010" , -- ADDR 206
			"00000000000011100110100010111000" , -- ADDR 207
			"00000000000000000110000110101000" , -- ADDR 208
			"00000000000001001011011111110001" , -- ADDR 209
			"00000000000010101010111010100111" , -- ADDR 210
			"00000000000001101001000110000001" , -- ADDR 211
			"00000000000001100001110110001100" , -- ADDR 212
			"00000000000001100011010001001010" , -- ADDR 213
			"00000000000010001100111010010010" , -- ADDR 214
			"00000000000001010001001010100101" , -- ADDR 215
			"00000000000001101010101001100011" , -- ADDR 216
			"00000000000000000111101110000111" , -- ADDR 217
			"00000000000000100100101001000011" , -- ADDR 218
			"00000000000010000110110101001100" , -- ADDR 219
			"00000000000010001110100111010001" , -- ADDR 220
			"00000000000001110100110110000000" , -- ADDR 221
			"00000000000001111100011100111011" , -- ADDR 222
			"00000000000010010001000110101100" , -- ADDR 223
			"00000000000001101010100101111110" , -- ADDR 224
			"00000000000001000001111101101001" , -- ADDR 225
			"00000000000010010000000010000110" , -- ADDR 226
			"00000000000000100111110110110000" , -- ADDR 227
			"00000000000000101001101110000000" , -- ADDR 228
			"00000000000000101000100101000000" , -- ADDR 229
			"00000000000000010101010110101000" , -- ADDR 230
			"00000000000000001100011100101110" , -- ADDR 231
			"00000000000000011110111001111110" , -- ADDR 232
			"00000000000000010100110010011011" , -- ADDR 233
			"00000000000001110101000100010001" , -- ADDR 234
			"00000000000011001110111100101011" , -- ADDR 235
			"00000000000001000001000111000101" , -- ADDR 236
			"00000000000000110011110100011010" , -- ADDR 237
			"00000000000001010000110111001010" , -- ADDR 238
			"00000000000000101001101010100100" , -- ADDR 239
			"00000000000010100100011100110111" , -- ADDR 240
			"00000000000000001011100101001010" , -- ADDR 241
			"00000000000000111011000011001100" , -- ADDR 242
			"00000000000001011110011001111101" , -- ADDR 243
			"00000000000001111010000011010101" , -- ADDR 244
			"00000000000011110000010101111001" , -- ADDR 245
			"00000000000011101001101001110000" , -- ADDR 246
			"00000000000001111000000000100010" , -- ADDR 247
			"00000000000010010001100000101000" , -- ADDR 248
			"00000000000001111111101111111011" , -- ADDR 249
			"00000000000010110001010001010111" , -- ADDR 250
			"00000000000001010101010001100101" , -- ADDR 251
			"00000000000010110101101100000010" , -- ADDR 252
			"00000000000011100001010010011101" , -- ADDR 253
			"00000000000000001001110101110111" , -- ADDR 254
			"00000000000001010000010001111000" , -- ADDR 255
			"00000000000010110011011100101001" , -- ADDR 256
			"00000000000001110001101100001000" , -- ADDR 257
			"00000000000001101000011110011011" , -- ADDR 258
			"00000000000001101010010000011110" , -- ADDR 259
			"00000000000010010101011000111111" , -- ADDR 260
			"00000000000001011001110001110010" , -- ADDR 261
			"00000000000001110010100001001100" , -- ADDR 262
			"00000000000000001101111010110001" , -- ADDR 263
			"00000000000000011110010100100101" , -- ADDR 264
			"00000000000010000010001101011011" , -- ADDR 265
			"00000000000010001000100000011001" , -- ADDR 266
			"00000000000001101110011001111001" , -- ADDR 267
			"00000000000010000000111010001111" , -- ADDR 268
			"00000000000010011000010001010011" , -- ADDR 269
			"00000000000001110011001100011000" , -- ADDR 270
			"00000000000001001010011110010001" , -- ADDR 271
			"00000000000010001010101110110011" , -- ADDR 272
			"00000000000000110000000101110001" , -- ADDR 273
			"00000000000000110010001011101100" , -- ADDR 274
			"00000000000000110001001001011100" , -- ADDR 275
			"00000000000000011101011111111110" , -- ADDR 276
			"00000000000000010101000100101001" , -- ADDR 277
			"00000000000000100111100010010101" , -- ADDR 278
			"00000000000000011101011001100000" , -- ADDR 279
			"00000000000001111011000011001001" , -- ADDR 280
			"00000000000011010111000110001100" , -- ADDR 281
			"00000000000000111111011111010000" , -- ADDR 282
			"00000000000000111010110011000000" , -- ADDR 283
			"00000000000001010111111010000101" , -- ADDR 284
			"00000000000000101100011011110011" , -- ADDR 285
			"00000000000010100001100110010110" , -- ADDR 286
			"00000000000000010001010000110111" , -- ADDR 287
			"00000000000001000011101011100010" , -- ADDR 288
			"00000000000001100101000001100001" , -- ADDR 289
			"00000000000001110001011010111010" , -- ADDR 290
			"00000000000011101001001000001111" , -- ADDR 291
			"00000000000011100000001001010000" , -- ADDR 292
			"00000000000100001011100011110100" , -- ADDR 293
			"00000000000100001011100000110010" , -- ADDR 294
			"00000000000110001101010100011101" , -- ADDR 295
			"00000000000100110000000000010001" , -- ADDR 296
			"00000000000101011111101000111000" , -- ADDR 297
			"00000000000101110011100000111110" , -- ADDR 298
			"00000000000011100100010111000001" , -- ADDR 299
			"00000000000010101110010010000111" , -- ADDR 300
			"00000000000001101110001010110000" , -- ADDR 301
			"00000000000010001001010001001010" , -- ADDR 302
			"00000000000011000101000001011001" , -- ADDR 303
			"00000000000010000110101101011010" , -- ADDR 304
			"00000000000001011000010100000100" , -- ADDR 305
			"00000000000010010100101101110011" , -- ADDR 306
			"00000000000001110111111010100100" , -- ADDR 307
			"00000000000011011100000000111100" , -- ADDR 308
			"00000000000011110111001011000111" , -- ADDR 309
			"00000000000100100010100011001111" , -- ADDR 310
			"00000000000100111100110101111011" , -- ADDR 311
			"00000000000100101101111100000100" , -- ADDR 312
			"00000000000010011011100000100101" , -- ADDR 313
			"00000000000001011110000111101111" , -- ADDR 314
			"00000000000001111100111000011101" , -- ADDR 315
			"00000000000010101011001100101111" , -- ADDR 316
			"00000000000101100100010110110000" , -- ADDR 317
			"00000000000010111001101000011001" , -- ADDR 318
			"00000000000010111000001000011101" , -- ADDR 319
			"00000000000010111001111011101001" , -- ADDR 320
			"00000000000011001100001011011100" , -- ADDR 321
			"00000000000011010101100011011010" , -- ADDR 322
			"00000000000011000100011000101010" , -- ADDR 323
			"00000000000011001110101011001001" , -- ADDR 324
			"00000000000011010001010111010011" , -- ADDR 325
			"00000000000000010010100101111110" , -- ADDR 326
			"00000000000100001011010010010110" , -- ADDR 327
			"00000000000010110001011111010101" , -- ADDR 328
			"00000000000011000000101110000111" , -- ADDR 329
			"00000000000011001110001010000111" , -- ADDR 330
			"00000000000100011010011011011100" , -- ADDR 331
			"00000000000011011001010101000111" , -- ADDR 332
			"00000000000010101011010100100010" , -- ADDR 333
			"00000000000010001110101110111101" , -- ADDR 334
			"00000000000101010111000010011000" , -- ADDR 335
			"00000000000110100010101101111010" , -- ADDR 336
			"00000000000000101100110010001111" , -- ADDR 337
			"00000000000000101100000001111011" , -- ADDR 338
			"00000000000100010111100001000110" , -- ADDR 339
			"00000000000011000110010000010010" , -- ADDR 340
			"00000000000100101101010110100110" , -- ADDR 341
			"00000000000101011001010001010111" , -- ADDR 342
			"00000000000001101110011111000100" , -- ADDR 343
			"00000000000010100001010111111000" , -- ADDR 344
			"00000000000001111011101011010110" , -- ADDR 345
			"00000000000001011101000100011111" , -- ADDR 346
			"00000000000000011110101111001001" , -- ADDR 347
			"00000000000010011011010000111100" , -- ADDR 348
			"00000000000010001101101100100100" , -- ADDR 349
			"00000000000001100101010100110110" , -- ADDR 350
			"00000000000010001111001111101000" , -- ADDR 351
			"00000000000001110110110010010000" , -- ADDR 352
			"00000000000010010110010001111101" , -- ADDR 353
			"00000000000011111001101101010011" , -- ADDR 354
			"00000000000100000000001100111101" , -- ADDR 355
			"00000000000011100101110000010101" , -- ADDR 356
			"00000000000011001010111000111111" , -- ADDR 357
			"00000000000010111001001111101101" , -- ADDR 358
			"00000000000001101111101000000100" , -- ADDR 359
			"00000000000001010010101100010111" , -- ADDR 360
			"00000000000010011101100000100011" , -- ADDR 361
			"00000000000001101111000101011000" , -- ADDR 362
			"00000000000001101010010100000100" , -- ADDR 363
			"00000000000001100110111010101001" , -- ADDR 364
			"00000000000001110000011100011010" , -- ADDR 365
			"00000000000001101100111000111010" , -- ADDR 366
			"00000000000001100101000010000000" , -- ADDR 367
			"00000000000001100110111011000110" , -- ADDR 368
			"00000000000000001111101000011111" , -- ADDR 369
			"00000000000011010000111100110110" , -- ADDR 370
			"00000000000001010111101001110010" , -- ADDR 371
			"00000000000010000001010101001101" , -- ADDR 372
			"00000000000000101101110000011001" , -- ADDR 373
			"00000000000010010010001000001100" , -- ADDR 374
			"00000000000100010101010100010100" , -- ADDR 375
			"00000000000001111000110111111101" , -- ADDR 376
			"00000000000001011101100111001110" , -- ADDR 377
			"00000000000010011101001011101001" , -- ADDR 378
			"00000000000011010001111111110001" , -- ADDR 379
			"00000000000101011101001111001000" , -- ADDR 380
			"00000000000000010100010100010001" , -- ADDR 381
			"00000000000100011100100100101011" , -- ADDR 382
			"00000000000011010101010110000000" , -- ADDR 383
			"00000000000101000001011110010101" , -- ADDR 384
			"00000000000101101111111100101100" , -- ADDR 385
			"00000000000010001001000100111111" , -- ADDR 386
			"00000000000011000111101100100011" , -- ADDR 387
			"00000000000010100011101001101101" , -- ADDR 388
			"00000000000010001001110110100110" , -- ADDR 389
			"00000000000001001011001101011010" , -- ADDR 390
			"00000000000011000101110100000111" , -- ADDR 391
			"00000000000010111010010101010001" , -- ADDR 392
			"00000000000010010000110010010011" , -- ADDR 393
			"00000000000010111011001001010111" , -- ADDR 394
			"00000000000010010100000000011110" , -- ADDR 395
			"00000000000010101110010111000010" , -- ADDR 396
			"00000000000100010010111011011111" , -- ADDR 397
			"00000000000100010100111111010100" , -- ADDR 398
			"00000000000011111010000111001111" , -- ADDR 399
			"00000000000011110011101101000011" , -- ADDR 400
			"00000000000011100101100111001100" , -- ADDR 401
			"00000000000010011100010100111000" , -- ADDR 402
			"00000000000001111100100001001001" , -- ADDR 403
			"00000000000010001011001101010101" , -- ADDR 404
			"00000000000010010100001100000100" , -- ADDR 405
			"00000000000010001111111001110100" , -- ADDR 406
			"00000000000010001100010011010010" , -- ADDR 407
			"00000000000010010001100001111011" , -- ADDR 408
			"00000000000010001011101000101100" , -- ADDR 409
			"00000000000010001000001100011101" , -- ADDR 410
			"00000000000010000111011111111000" , -- ADDR 411
			"00000000000000111010011010100110" , -- ADDR 412
			"00000000000011111100110101001000" , -- ADDR 413
			"00000000000001011111001100110000" , -- ADDR 414
			"00000000000010100111011000010000" , -- ADDR 415
			"00000000000001011000000110100011" , -- ADDR 416
			"00000000000010110011001011000110" , -- ADDR 417
			"00000000000100110010111001100100" , -- ADDR 418
			"00000000000010010110110101101111" , -- ADDR 419
			"00000000000010000110011010101000" , -- ADDR 420
			"00000000000011000111000000100010" , -- ADDR 421
			"00000000000011010111101000100001" , -- ADDR 422
			"00000000000101101010111110110111" , -- ADDR 423
			"00000000000100001000010100010111" , -- ADDR 424
			"00000000000011000001011000010110" , -- ADDR 425
			"00000000000100101101111001100010" , -- ADDR 426
			"00000000000101011100101101000110" , -- ADDR 427
			"00000000000001110111101111000001" , -- ADDR 428
			"00000000000010111010011100101100" , -- ADDR 429
			"00000000000010100111100110001101" , -- ADDR 430
			"00000000000010000101110001101111" , -- ADDR 431
			"00000000000001000111000001011000" , -- ADDR 432
			"00000000000010111100000011100100" , -- ADDR 433
			"00000000000010110111011101111010" , -- ADDR 434
			"00000000000010001000110010100010" , -- ADDR 435
			"00000000000010110011011011010100" , -- ADDR 436
			"00000000000010000011010011011100" , -- ADDR 437
			"00000000000010011011111101111111" , -- ADDR 438
			"00000000000100000000010101111000" , -- ADDR 439
			"00000000000100000001100101000111" , -- ADDR 440
			"00000000000011100110101100100110" , -- ADDR 441
			"00000000000011100111111100100101" , -- ADDR 442
			"00000000000011011110101100001100" , -- ADDR 443
			"00000000000010010111001100011110" , -- ADDR 444
			"00000000000001110010111111100010" , -- ADDR 445
			"00000000000001111010010010100011" , -- ADDR 446
			"00000000000010000110110101001100" , -- ADDR 447
			"00000000000010000010111001010000" , -- ADDR 448
			"00000000000001111111001111011001" , -- ADDR 449
			"00000000000010000010010010100011" , -- ADDR 450
			"00000000000001111011100101100011" , -- ADDR 451
			"00000000000001111010000011010101" , -- ADDR 452
			"00000000000001111000001110011011" , -- ADDR 453
			"00000000000000111011100100001001" , -- ADDR 454
			"00000000000011111011111100010000" , -- ADDR 455
			"00000000000001001011001000111110" , -- ADDR 456
			"00000000000010011010010010101101" , -- ADDR 457
			"00000000000001010000010100110110" , -- ADDR 458
			"00000000000010100011011111001101" , -- ADDR 459
			"00000000000100100001010110010001" , -- ADDR 460
			"00000000000010000110010110000001" , -- ADDR 461
			"00000000000001111011110001111001" , -- ADDR 462
			"00000000000010111100011101111010" , -- ADDR 463
			"00000000000011000011010101001110" , -- ADDR 464
			"00000000000101010110110010000111" , -- ADDR 465
			"00000000000001011110100000000000" , -- ADDR 466
			"00000000000001101100000101011111" , -- ADDR 467
			"00000000000010010111010000100100" , -- ADDR 468
			"00000000000010111010000111111101" , -- ADDR 469
			"00000000000011011111010110000110" , -- ADDR 470
			"00000000000101100100100111010101" , -- ADDR 471
			"00000000000100100010100011001111" , -- ADDR 472
			"00000000000100010010011111001100" , -- ADDR 473
			"00000000000100000110100111001111" , -- ADDR 474
			"00000000000101000000110101111101" , -- ADDR 475
			"00000000000100001001000001111100" , -- ADDR 476
			"00000000000100010111001011100101" , -- ADDR 477
			"00000000000010111011111111100000" , -- ADDR 478
			"00000000000010011010000111100101" , -- ADDR 479
			"00000000000010000100000101110001" , -- ADDR 480
			"00000000000001100101111010011001" , -- ADDR 481
			"00000000000001100101111101101010" , -- ADDR 482
			"00000000000011111110011111101101" , -- ADDR 483
			"00000000000100110001011010011010" , -- ADDR 484
			"00000000000100100001101111011101" , -- ADDR 485
			"00000000000011111011101101000111" , -- ADDR 486
			"00000000000010101100011001010110" , -- ADDR 487
			"00000000000011011101001010011100" , -- ADDR 488
			"00000000000011100000101100010100" , -- ADDR 489
			"00000000000011100000100111110110" , -- ADDR 490
			"00000000000011001011110111110100" , -- ADDR 491
			"00000000000011000101110110010010" , -- ADDR 492
			"00000000000011011000000110000111" , -- ADDR 493
			"00000000000011001110011011011100" , -- ADDR 494
			"00000000000100100000000110001010" , -- ADDR 495
			"00000000000101111010111111000001" , -- ADDR 496
			"00000000000011000000101011111000" , -- ADDR 497
			"00000000000011011110111000011001" , -- ADDR 498
			"00000000000100000100101110110010" , -- ADDR 499
			"00000000000011000000000011101110" , -- ADDR 500
			"00000000000010101100001010001000" , -- ADDR 501
			"00000000000010111101001110011001" , -- ADDR 502
			"00000000000011110100001001001100" , -- ADDR 503
			"00000000000011111110100111110001" , -- ADDR 504
			"00000000000001000101100101110100" , -- ADDR 505
			"00000000000001100001010011100000" , -- ADDR 506
			"00000000000001101110011000100110" , -- ADDR 507
			"00000000000010011111011110111010" , -- ADDR 508
			"00000000000001011110110000001000" , -- ADDR 509
			"00000000000010000011010001100111" , -- ADDR 510
			"00000000000100000111010001010011" , -- ADDR 511
			"00000000000011000100111111011101" , -- ADDR 512
			"00000000000010111011101101001111" , -- ADDR 513
			"00000000000010101001011101111000" , -- ADDR 514
			"00000000000011100010010110111000" , -- ADDR 515
			"00000000000010101010111001110010" , -- ADDR 516
			"00000000000010111001000110011100" , -- ADDR 517
			"00000000000001011110101000100101" , -- ADDR 518
			"00000000000000111011110100001000" , -- ADDR 519
			"00000000000001010001110010111101" , -- ADDR 520
			"00000000000001000101001001101000" , -- ADDR 521
			"00000000000000101100100011010011" , -- ADDR 522
			"00000000000010101000000000111010" , -- ADDR 523
			"00000000000011010101100010010011" , -- ADDR 524
			"00000000000011000011011010000111" , -- ADDR 525
			"00000000000010011110110101010001" , -- ADDR 526
			"00000000000010001110101000010001" , -- ADDR 527
			"00000000000001111110111101000000" , -- ADDR 528
			"00000000000010000010101010101010" , -- ADDR 529
			"00000000000010000010110100100000" , -- ADDR 530
			"00000000000001101110000110110111" , -- ADDR 531
			"00000000000001101000111101110110" , -- ADDR 532
			"00000000000001111010110011101000" , -- ADDR 533
			"00000000000001110001100110010000" , -- ADDR 534
			"00000000000011001100001011011100" , -- ADDR 535
			"00000000000100011101100011011010" , -- ADDR 536
			"00000000000001110110010000011101" , -- ADDR 537
			"00000000000010000000011100100110" , -- ADDR 538
			"00000000000010101100001100010101" , -- ADDR 539
			"00000000000001100001111111111100" , -- ADDR 540
			"00000000000001111110010100101101" , -- ADDR 541
			"00000000000001011111011111110000" , -- ADDR 542
			"00000000000010010110100011000100" , -- ADDR 543
			"00000000000010100001110000111110" , -- ADDR 544
			"00000000000000101101111100110111" , -- ADDR 545
			"00000000000010010111000001000111" , -- ADDR 546
			"00000000000000110010001011101100" , -- ADDR 547
			"00000000000010111111011011011100" , -- ADDR 548
			"00000000000010111001010111101100" , -- ADDR 549
			"00000000000101010101101011010101" , -- ADDR 550
			"00000000000100010101011110011101" , -- ADDR 551
			"00000000000100011101100000111010" , -- ADDR 552
			"00000000000011100000100101101110" , -- ADDR 553
			"00000000000100100011101100000111" , -- ADDR 554
			"00000000000011111001001000000001" , -- ADDR 555
			"00000000000011110110001000111111" , -- ADDR 556
			"00000000000010111001100010001111" , -- ADDR 557
			"00000000000010010111011000110001" , -- ADDR 558
			"00000000000000111110000001000010" , -- ADDR 559
			"00000000000000101101001011101100" , -- ADDR 560
			"00000000000001000111101100001001" , -- ADDR 561
			"00000000000011000100100110000000" , -- ADDR 562
			"00000000000100000001110110111000" , -- ADDR 563
			"00000000000100001101011100100101" , -- ADDR 564
			"00000000000011110101001001111010" , -- ADDR 565
			"00000000000011110110101010110111" , -- ADDR 566
			"00000000000011010000100010100101" , -- ADDR 567
			"00000000000011010101011101001010" , -- ADDR 568
			"00000000000011010111001000101000" , -- ADDR 569
			"00000000000011000101000000001011" , -- ADDR 570
			"00000000000011000100010111011100" , -- ADDR 571
			"00000000000011010010100111101011" , -- ADDR 572
			"00000000000011001100001100011000" , -- ADDR 573
			"00000000000100110000101101001111" , -- ADDR 574
			"00000000000101001110110010110001" , -- ADDR 575
			"00000000000011100011010000101100" , -- ADDR 576
			"00000000000011001000100111011001" , -- ADDR 577
			"00000000000100001100001001011000" , -- ADDR 578
			"00000000000010101001111011011000" , -- ADDR 579
			"00000000000001001111001101000111" , -- ADDR 580
			"00000000000010111000100010010100" , -- ADDR 581
			"00000000000011101010001100110100" , -- ADDR 582
			"00000000000011010111111101101110" , -- ADDR 583
			"00000000000010000011110000011100" , -- ADDR 584
			"00000000000001000100000010000001" , -- ADDR 585
			"00000000000011101010110010011011" , -- ADDR 586
			"00000000000011010111110010101011" , -- ADDR 587
			"00000000000101110110100100001010" , -- ADDR 588
			"00000000000100111000101010100010" , -- ADDR 589
			"00000000000101000111010011011010" , -- ADDR 590
			"00000000000011111100100110011010" , -- ADDR 591
			"00000000000101000000100110110010" , -- ADDR 592
			"00000000000100011100010110010001" , -- ADDR 593
			"00000000000100010011001100101001" , -- ADDR 594
			"00000000000011100011011000011101" , -- ADDR 595
			"00000000000011000011000110110100" , -- ADDR 596
			"00000000000001100000101011101011" , -- ADDR 597
			"00000000000001011011011010100001" , -- ADDR 598
			"00000000000001110110001101001111" , -- ADDR 599
			"00000000000011011000101010000010" , -- ADDR 600
			"00000000000100010111111001110100" , -- ADDR 601
			"00000000000100101110011100000110" , -- ADDR 602
			"00000000000100011011011010101001" , -- ADDR 603
			"00000000000100101000110110100001" , -- ADDR 604
			"00000000000011110110100000110011" , -- ADDR 605
			"00000000000011111011100111000010" , -- ADDR 606
			"00000000000011111101101110010111" , -- ADDR 607
			"00000000000011101101001010001100" , -- ADDR 608
			"00000000000011101101111011111110" , -- ADDR 609
			"00000000000011111010100001101110" , -- ADDR 610
			"00000000000011110101001110100101" , -- ADDR 611
			"00000000000101011011011011000011" , -- ADDR 612
			"00000000000101100011110101001001" , -- ADDR 613
			"00000000000100010010101110011110" , -- ADDR 614
			"00000000000011101011111011111110" , -- ADDR 615
			"00000000000100110101011101101111" , -- ADDR 616
			"00000000000011001111001101111100" , -- ADDR 617
			"00000000000001011001000110100110" , -- ADDR 618
			"00000000000011100001111000100000" , -- ADDR 619
			"00000000000100001111110111011100" , -- ADDR 620
			"00000000000011110100001010111101" , -- ADDR 621
			"00000000000010110101110011001000" , -- ADDR 622
			"00000000000001001101110110111000" , -- ADDR 623
			"00000000000001010001001001111111" , -- ADDR 624
			"00000000000010101010111100000001" , -- ADDR 625
			"00000000000001101001100011011100" , -- ADDR 626
			"00000000000001011110101000100101" , -- ADDR 627
			"00000000000001100111101101011010" , -- ADDR 628
			"00000000000010001111000010010011" , -- ADDR 629
			"00000000000001010010101010101000" , -- ADDR 630
			"00000000000001101110000111101110" , -- ADDR 631
			"00000000000000001101101001011110" , -- ADDR 632
			"00000000000000101000000010101100" , -- ADDR 633
			"00000000000010001011011011000010" , -- ADDR 634
			"00000000000010010010010000000001" , -- ADDR 635
			"00000000000001111000001101001111" , -- ADDR 636
			"00000000000010000010001010001000" , -- ADDR 637
			"00000000000010010101010101001010" , -- ADDR 638
			"00000000000001101100001001111001" , -- ADDR 639
			"00000000000001000010000001010000" , -- ADDR 640
			"00000000000010001010110110000001" , -- ADDR 641
			"00000000000000101011000000001011" , -- ADDR 642
			"00000000000000101100001110111001" , -- ADDR 643
			"00000000000000101010101000110010" , -- ADDR 644
			"00000000000000011001000010111111" , -- ADDR 645
			"00000000000000001110111001101001" , -- ADDR 646
			"00000000000000100000011011110101" , -- ADDR 647
			"00000000000000010110000000011011" , -- ADDR 648
			"00000000000001110001010010000100" , -- ADDR 649
			"00000000000011010001110111001001" , -- ADDR 650
			"00000000000000111011000011001100" , -- ADDR 651
			"00000000000000111000011011100010" , -- ADDR 652
			"00000000000001001110000110001011" , -- ADDR 653
			"00000000000000101111101111111000" , -- ADDR 654
			"00000000000010101001110100101001" , -- ADDR 655
			"00000000000000010001011110100101" , -- ADDR 656
			"00000000000000111100000111001101" , -- ADDR 657
			"00000000000001100011001000111111" , -- ADDR 658
			"00000000000001111001010110010001" , -- ADDR 659
			"00000000000011110010111100101001" , -- ADDR 660
			"00000000000010011110110111010111" , -- ADDR 661
			"00000000000001100011100100010110" , -- ADDR 662
			"00000000000010000101111111111110" , -- ADDR 663
			"00000000000000101000010011010100" , -- ADDR 664
			"00000000000001101010010100100000" , -- ADDR 665
			"00000000000001001000100001101101" , -- ADDR 666
			"00000000000000111100110100001010" , -- ADDR 667
			"00000000000001000011110011010010" , -- ADDR 668
			"00000000000001001111101101100001" , -- ADDR 669
			"00000000000001111011011101011101" , -- ADDR 670
			"00000000000010010001111000100001" , -- ADDR 671
			"00000000000010000000011000100000" , -- ADDR 672
			"00000000000000110001000001101011" , -- ADDR 673
			"00000000000001010010010010111011" , -- ADDR 674
			"00000000000001010111000101110001" , -- ADDR 675
			"00000000000001010000110011000010" , -- ADDR 676
			"00000000000011011011000000101001" , -- ADDR 677
			"00000000000000110011101000011011" , -- ADDR 678
			"00000000000000110111110010110000" , -- ADDR 679
			"00000000000000111011011001101111" , -- ADDR 680
			"00000000000000111011100111010110" , -- ADDR 681
			"00000000000001000101010001111001" , -- ADDR 682
			"00000000000001000000101101010111" , -- ADDR 683
			"00000000000001000100111001000011" , -- ADDR 684
			"00000000000010011100011100001101" , -- ADDR 685
			"00000000000010011100001000101011" , -- ADDR 686
			"00000000000010001011001011101000" , -- ADDR 687
			"00000000000000100000010100011110" , -- ADDR 688
			"00000000000001110100010011001110" , -- ADDR 689
			"00000000000000100110000001001100" , -- ADDR 690
			"00000000000010000011101101100011" , -- ADDR 691
			"00000000000000111111111101001100" , -- ADDR 692
			"00000000000001000100110011100000" , -- ADDR 693
			"00000000000000011111110101010000" , -- ADDR 694
			"00000000000010101101010111011010" , -- ADDR 695
			"00000000000011111001101011001100" , -- ADDR 696
			"00000000000001000010010100101110" , -- ADDR 697
			"00000000000001100110110011101100" , -- ADDR 698
			"00000000000001111101000001001111" , -- ADDR 699
			"00000000000000111101110001101000" , -- ADDR 700
			"00000000000001011101100111001110" , -- ADDR 701
			"00000000000001100110000011010001" , -- ADDR 702
			"00000000000010101000101111010110" , -- ADDR 703
			"00000000000011001011101100100101" , -- ADDR 704
			"00000000000100011000101000100110" , -- ADDR 705
			"00000000000100101011010100100100" , -- ADDR 706
			"00000000000100010101011011001100" , -- ADDR 707
			"00000000000010101100101101100001" , -- ADDR 708
			"00000000000001111000001101101000" , -- ADDR 709
			"00000000000001001000010011111000" , -- ADDR 710
			"00000000000001101000111110110000" , -- ADDR 711
			"00000000000100010001100000100010" , -- ADDR 712
			"00000000000010001001000100111111" , -- ADDR 713
			"00000000000010000100111100000110" , -- ADDR 714
			"00000000000010000100100001001010" , -- ADDR 715
			"00000000000010011001001011010111" , -- ADDR 716
			"00000000000010011110110001000100" , -- ADDR 717
			"00000000000010001100100100100110" , -- ADDR 718
			"00000000000010010110001100001111" , -- ADDR 719
			"00000000000001101100000100001010" , -- ADDR 720
			"00000000000001100011101000001011" , -- ADDR 721
			"00000000000010111100110010001000" , -- ADDR 722
			"00000000000010001101010111000000" , -- ADDR 723
			"00000000000001101010100101100010" , -- ADDR 724
			"00000000000010101100111010011111" , -- ADDR 725
			"00000000000100100001111101110001" , -- ADDR 726
			"00000000000010100111110001100100" , -- ADDR 727
			"00000000000001110000101110101000" , -- ADDR 728
			"00000000000010000100101110000110" , -- ADDR 729
			"00000000000100100100000111011001" , -- ADDR 730
			"00000000000110010010101011011011" , -- ADDR 731
			"00000000000000111111000001000110" , -- ADDR 732
			"00000000000001001010110100101000" , -- ADDR 733
			"00000000000000110010000110111100" , -- ADDR 734
			"00000000000000011100011001001001" , -- ADDR 735
			"00000000000000111000000000011001" , -- ADDR 736
			"00000000000001100110100100010111" , -- ADDR 737
			"00000000000010001001011000000110" , -- ADDR 738
			"00000000000011011001010010010000" , -- ADDR 739
			"00000000000011101010010110100101" , -- ADDR 740
			"00000000000011010011110001101111" , -- ADDR 741
			"00000000000001111110001010100001" , -- ADDR 742
			"00000000000001011110000000001000" , -- ADDR 743
			"00000000000000010011100100011100" , -- ADDR 744
			"00000000000000100111101111100100" , -- ADDR 745
			"00000000000011011100100001001100" , -- ADDR 746
			"00000000000001000110110111010011" , -- ADDR 747
			"00000000000001000010101000110011" , -- ADDR 748
			"00000000000001000010001100110011" , -- ADDR 749
			"00000000000001010110111000100111" , -- ADDR 750
			"00000000000001011100110011100100" , -- ADDR 751
			"00000000000001001010011101101000" , -- ADDR 752
			"00000000000001010100010011101110" , -- ADDR 753
			"00000000000001010000101011111100" , -- ADDR 754
			"00000000000001111000010110110000" , -- ADDR 755
			"00000000000010000100000111001101" , -- ADDR 756
			"00000000000001001100111111011101" , -- ADDR 757
			"00000000000000110111101011000011" , -- ADDR 758
			"00000000000001101011101110111101" , -- ADDR 759
			"00000000000011100110111101010101" , -- ADDR 760
			"00000000000001100101100000001000" , -- ADDR 761
			"00000000000000101110011100110111" , -- ADDR 762
			"00000000000001010000001111100000" , -- ADDR 763
			"00000000000011100010111001011000" , -- ADDR 764
			"00000000000101010001001101010100" , -- ADDR 765
			"00000000000001111101000110111101" , -- ADDR 766
			"00000000000001110000011101101100" , -- ADDR 767
			"00000000000001000110110101111100" , -- ADDR 768
			"00000000000001110000100010110001" , -- ADDR 769
			"00000000000001100100000110101110" , -- ADDR 770
			"00000000000010000110011100011001" , -- ADDR 771
			"00000000000011100110110101000100" , -- ADDR 772
			"00000000000011110000011010011101" , -- ADDR 773
			"00000000000011010110101011100100" , -- ADDR 774
			"00000000000010101101100101011011" , -- ADDR 775
			"00000000000010011010100001110101" , -- ADDR 776
			"00000000000001010001001001111111" , -- ADDR 777
			"00000000000000110101101010110101" , -- ADDR 778
			"00000000000010101011000010101101" , -- ADDR 779
			"00000000000001010101101010101100" , -- ADDR 780
			"00000000000001010000100111001101" , -- ADDR 781
			"00000000000001001101100010000001" , -- ADDR 782
			"00000000000001011010101000110000" , -- ADDR 783
			"00000000000001011001011010010111" , -- ADDR 784
			"00000000000001001101110110111000" , -- ADDR 785
			"00000000000001010010000111010101" , -- ADDR 786
			"00000000000000010110011100010100" , -- ADDR 787
			"00000000000010110101001000100011" , -- ADDR 788
			"00000000000001011001110010010100" , -- ADDR 789
			"00000000000001100110101000100011" , -- ADDR 790
			"00000000000000010010010011111000" , -- ADDR 791
			"00000000000001111011001010100000" , -- ADDR 792
			"00000000000011111111000101101100" , -- ADDR 793
			"00000000000001100101011011111010" , -- ADDR 794
			"00000000000001000001010010110010" , -- ADDR 795
			"00000000000001111111011011101111" , -- ADDR 796
			"00000000000011001101111010110101" , -- ADDR 797
			"00000000000101010001011001000011" , -- ADDR 798
			"00000000000001000100000000101000" , -- ADDR 799
			"00000000000000110110100101110111" , -- ADDR 800
			"00000000000000010111000010000100" , -- ADDR 801
			"00000000000001011100011001010011" , -- ADDR 802
			"00000000000001110010000110111010" , -- ADDR 803
			"00000000000010100010100100101110" , -- ADDR 804
			"00000000000010111001111100101011" , -- ADDR 805
			"00000000000010101000101011000111" , -- ADDR 806
			"00000000000000110011010101111001" , -- ADDR 807
			"00000000000000101110001001010011" , -- ADDR 808
			"00000000000000111001100111101000" , -- ADDR 809
			"00000000000001001001010101010111" , -- ADDR 810
			"00000000000011110001101100111101" , -- ADDR 811
			"00000000000000111110101000110100" , -- ADDR 812
			"00000000000000111111111010001101" , -- ADDR 813
			"00000000000001000011001001100101" , -- ADDR 814
			"00000000000001001110110001111100" , -- ADDR 815
			"00000000000001011001001111101100" , -- ADDR 816
			"00000000000001001100100111110111" , -- ADDR 817
			"00000000000001010101000000001110" , -- ADDR 818
			"00000000000010010010101111010001" , -- ADDR 819
			"00000000000001110100011000100011" , -- ADDR 820
			"00000000000010011011110011010001" , -- ADDR 821
			"00000000000000101111011110110111" , -- ADDR 822
			"00000000000001101101110111101100" , -- ADDR 823
			"00000000000001001000001000101010" , -- ADDR 824
			"00000000000010100101111101100011" , -- ADDR 825
			"00000000000001011001000000101101" , -- ADDR 826
			"00000000000001000000011010111001" , -- ADDR 827
			"00000000000000001000101000011011" , -- ADDR 828
			"00000000000011010001101110111101" , -- ADDR 829
			"00000000000100100001100100100110" , -- ADDR 830
			"00000000000000111101001011100111" , -- ADDR 831
			"00000000000000101101100110111111" , -- ADDR 832
			"00000000000010001000010101001101" , -- ADDR 833
			"00000000000010100111001010110110" , -- ADDR 834
			"00000000000011100101110000010101" , -- ADDR 835
			"00000000000011111011101100111010" , -- ADDR 836
			"00000000000011101000011110011101" , -- ADDR 837
			"00000000000001110000000110010101" , -- ADDR 838
			"00000000000000111010111101100010" , -- ADDR 839
			"00000000000000100100100111110000" , -- ADDR 840
			"00000000000001010011000001000101" , -- ADDR 841
			"00000000000100001100000011101100" , -- ADDR 842
			"00000000000001100101100111001011" , -- ADDR 843
			"00000000000001100011001101010100" , -- ADDR 844
			"00000000000001100100011100001000" , -- ADDR 845
			"00000000000001111000000101010011" , -- ADDR 846
			"00000000000010000000100101110111" , -- ADDR 847
			"00000000000001101110100111101100" , -- ADDR 848
			"00000000000001111001000010111111" , -- ADDR 849
			"00000000000010000000001011100000" , -- ADDR 850
			"00000000000001000110110001111010" , -- ADDR 851
			"00000000000010110011000000111110" , -- ADDR 852
			"00000000000001100010000001111000" , -- ADDR 853
			"00000000000001101001101110010010" , -- ADDR 854
			"00000000000010000001011111001001" , -- ADDR 855
			"00000000000011101001110001101101" , -- ADDR 856
			"00000000000010000110001001100101" , -- ADDR 857
			"00000000000001010100000101100100" , -- ADDR 858
			"00000000000001001100011100101001" , -- ADDR 859
			"00000000000100000101101110000111" , -- ADDR 860
			"00000000000101100011101001000101" , -- ADDR 861
			"00000000000000101010101000110010" , -- ADDR 862
			"00000000000001001101100001011010" , -- ADDR 863
			"00000000000001101111000101110011" , -- ADDR 864
			"00000000000010111100111001001101" , -- ADDR 865
			"00000000000011001110001000101110" , -- ADDR 866
			"00000000000010110111110110110101" , -- ADDR 867
			"00000000000001101000100111100011" , -- ADDR 868
			"00000000000001010110000101010110" , -- ADDR 869
			"00000000000000011001011111010011" , -- ADDR 870
			"00000000000000010111101100111010" , -- ADDR 871
			"00000000000011010000001111010111" , -- ADDR 872
			"00000000000000101011111101100101" , -- ADDR 873
			"00000000000000101000010110110111" , -- ADDR 874
			"00000000000000101000101111100011" , -- ADDR 875
			"00000000000000111101010101101111" , -- ADDR 876
			"00000000000001000100101101111101" , -- ADDR 877
			"00000000000000110010010101001011" , -- ADDR 878
			"00000000000000111100101101000110" , -- ADDR 879
			"00000000000001011100001101011010" , -- ADDR 880
			"00000000000010000010100111101111" , -- ADDR 881
			"00000000000001110111001010101101" , -- ADDR 882
			"00000000000000110000100110010100" , -- ADDR 883
			"00000000000000111000110011001000" , -- ADDR 884
			"00000000000001001111100001100010" , -- ADDR 885
			"00000000000011001011001110010110" , -- ADDR 886
			"00000000000001001011111011011110" , -- ADDR 887
			"00000000000000010110111011110101" , -- ADDR 888
			"00000000000000111001111001110011" , -- ADDR 889
			"00000000000011001011000101111001" , -- ADDR 890
			"00000000000100110101001100111011" , -- ADDR 891
			"00000000000001100100101100101110" , -- ADDR 892
			"00000000000001111111011000110000" , -- ADDR 893
			"00000000000010111000001011100100" , -- ADDR 894
			"00000000000011001110100001101011" , -- ADDR 895
			"00000000000010111100000001100010" , -- ADDR 896
			"00000000000001001000010001001111" , -- ADDR 897
			"00000000000000101011110000100010" , -- ADDR 898
			"00000000000000100101001011111011" , -- ADDR 899
			"00000000000001000001010010110010" , -- ADDR 900
			"00000000000011110100100111101001" , -- ADDR 901
			"00000000000001000011001000111000" , -- ADDR 902
			"00000000000001000010100110101001" , -- ADDR 903
			"00000000000001000101000100110011" , -- ADDR 904
			"00000000000001010101010100011000" , -- ADDR 905
			"00000000000001011111001110010000" , -- ADDR 906
			"00000000000001001111011111001000" , -- ADDR 907
			"00000000000001011001001111101100" , -- ADDR 908
			"00000000000010000101000011111111" , -- ADDR 909
			"00000000000001100101010100110110" , -- ADDR 910
			"00000000000010011100100001101100" , -- ADDR 911
			"00000000000000111001100101001010" , -- ADDR 912
			"00000000000001100011010110111011" , -- ADDR 913
			"00000000000001010111001001000011" , -- ADDR 914
			"00000000000010111100111000111100" , -- ADDR 915
			"00000000000001100001110100010000" , -- ADDR 916
			"00000000000000111011101010100011" , -- ADDR 917
			"00000000000000011111000111110011" , -- ADDR 918
			"00000000000011011111001011110110" , -- ADDR 919
			"00000000000100110110011001111001" , -- ADDR 920
			"00000000000000100011111001101110" , -- ADDR 921
			"00000000000010000011001100111001" , -- ADDR 922
			"00000000000010001100100001111000" , -- ADDR 923
			"00000000000001110011010000000110" , -- ADDR 924
			"00000000000001110100101111011110" , -- ADDR 925
			"00000000000010001010011000000101" , -- ADDR 926
			"00000000000001100110101111111110" , -- ADDR 927
			"00000000000001000000001110010011" , -- ADDR 928
			"00000000000010010111100100101110" , -- ADDR 929
			"00000000000000100010101111011110" , -- ADDR 930
			"00000000000000100101010110001011" , -- ADDR 931
			"00000000000000100100110011011100" , -- ADDR 932
			"00000000000000010000010010010100" , -- ADDR 933
			"00000000000000001010111010110001" , -- ADDR 934
			"00000000000000011100001011101010" , -- ADDR 935
			"00000000000000010011010011010001" , -- ADDR 936
			"00000000000001111000000011101101" , -- ADDR 937
			"00000000000011001001011100100001" , -- ADDR 938
			"00000000000001001000101011100100" , -- ADDR 939
			"00000000000000101100111010110000" , -- ADDR 940
			"00000000000001010010100111001010" , -- ADDR 941
			"00000000000000100010001100111001" , -- ADDR 942
			"00000000000010011111010100001001" , -- ADDR 943
			"00000000000000000011110111000011" , -- ADDR 944
			"00000000000000111000001001110000" , -- ADDR 945
			"00000000000001010111010010010110" , -- ADDR 946
			"00000000000001111101101011110110" , -- ADDR 947
			"00000000000011101111101000100110" , -- ADDR 948
			"00000000000001100100100111000010" , -- ADDR 949
			"00000000000001101010001101010101" , -- ADDR 950
			"00000000000001010000001111100000" , -- ADDR 951
			"00000000000001111100010011010101" , -- ADDR 952
			"00000000000010011111101111101001" , -- ADDR 953
			"00000000000010000111101000101011" , -- ADDR 954
			"00000000000001100011110101100100" , -- ADDR 955
			"00000000000010010011111010000010" , -- ADDR 956
			"00000000000001000011001000111000" , -- ADDR 957
			"00000000000001000110111001010100" , -- ADDR 958
			"00000000000001000111001011011100" , -- ADDR 959
			"00000000000000110010100101001111" , -- ADDR 960
			"00000000000000101110101110010001" , -- ADDR 961
			"00000000000000111111101100000000" , -- ADDR 962
			"00000000000000110111001100111100" , -- ADDR 963
			"00000000000010011001010100101101" , -- ADDR 964
			"00000000000011100100100110111000" , -- ADDR 965
			"00000000000001010110100001100001" , -- ADDR 966
			"00000000000001000101111011000000" , -- ADDR 967
			"00000000000001110101011111111010" , -- ADDR 968
			"00000000000000101010010100100101" , -- ADDR 969
			"00000000000010000110011100011001" , -- ADDR 970
			"00000000000000100100001001100111" , -- ADDR 971
			"00000000000001011010111111110110" , -- ADDR 972
			"00000000000001101011001100110010" , -- ADDR 973
			"00000000000001011111111000101011" , -- ADDR 974
			"00000000000011001011111000111111" , -- ADDR 975
			"00000000000000011110110011110010" , -- ADDR 976
			"00000000000000100110110010110110" , -- ADDR 977
			"00000000000010001000011011001001" , -- ADDR 978
			"00000000000011000100100010011000" , -- ADDR 979
			"00000000000011010000010100110110" , -- ADDR 980
			"00000000000010111010111001000010" , -- ADDR 981
			"00000000000011011111111100111010" , -- ADDR 982
			"00000000000010010101111111100010" , -- ADDR 983
			"00000000000010011011000100000010" , -- ADDR 984
			"00000000000010011101000111000101" , -- ADDR 985
			"00000000000010001100100000110111" , -- ADDR 986
			"00000000000010001101100110100000" , -- ADDR 987
			"00000000000010011001110110100011" , -- ADDR 988
			"00000000000010010100101101110011" , -- ADDR 989
			"00000000000011111011001110000000" , -- ADDR 990
			"00000000000100010001011101100100" , -- ADDR 991
			"00000000000010111000100001010010" , -- ADDR 992
			"00000000000010001100010011010010" , -- ADDR 993
			"00000000000011010100111010000011" , -- ADDR 994
			"00000000000001101110110000101111" , -- ADDR 995
			"00000000000000101101010011000100" , -- ADDR 996
			"00000000000010000001100001010111" , -- ADDR 997
			"00000000000010101111011101010111" , -- ADDR 998
			"00000000000010011001111100101111" , -- ADDR 999
			"00000000000001111001000110001001" , -- ADDR 1000
			"00000000000010000000001011001000" , -- ADDR 1001
			"00000000000000011010111000100010" , -- ADDR 1002
			"00000000000010100100011110000001" , -- ADDR 1003
			"00000000000011011110101110111110" , -- ADDR 1004
			"00000000000011100011011001111010" , -- ADDR 1005
			"00000000000011001000111101001111" , -- ADDR 1006
			"00000000000011010010011011101011" , -- ADDR 1007
			"00000000000010100100100111010011" , -- ADDR 1008
			"00000000000010101001011011101000" , -- ADDR 1009
			"00000000000010101010111100010011" , -- ADDR 1010
			"00000000000010011000010111110111" , -- ADDR 1011
			"00000000000010010111011001000101" , -- ADDR 1012
			"00000000000010100110000001000000" , -- ADDR 1013
			"00000000000010011111010100001001" , -- ADDR 1014
			"00000000000100000011100001111110" , -- ADDR 1015
			"00000000000100101011010111111010" , -- ADDR 1016
			"00000000000010110111010110111001" , -- ADDR 1017
			"00000000000010011101111101100100" , -- ADDR 1018
			"00000000000011011111000111110010" , -- ADDR 1019
			"00000000000001111110100111111100" , -- ADDR 1020
			"00000000000001000111001011011100" , -- ADDR 1021
			"00000000000010001011101000101100" , -- ADDR 1022
			"00000000000010111110010000101111" , -- ADDR 1023
			"00000000000010110001010101111011" , -- ADDR 1024
			"00000000000001100100001101111000" , -- ADDR 1025
			"00000000000001100111111101000001" , -- ADDR 1026
			"00000000000010011001101110110010" , -- ADDR 1027
			"00000000000011010000010100101000" , -- ADDR 1028
			"00000000000011001110001000111101" , -- ADDR 1029
			"00000000000010110001000010100011" , -- ADDR 1030
			"00000000000010111011001001010111" , -- ADDR 1031
			"00000000000010001101010010010001" , -- ADDR 1032
			"00000000000010010001111011001000" , -- ADDR 1033
			"00000000000010010011001010001100" , -- ADDR 1034
			"00000000000001111111111010010111" , -- ADDR 1035
			"00000000000001111110001010100001" , -- ADDR 1036
			"00000000000010001101100010110011" , -- ADDR 1037
			"00000000000010000110010011001011" , -- ADDR 1038
			"00000000000011101001011011110111" , -- ADDR 1039
			"00000000000100011100000010111110" , -- ADDR 1040
			"00000000000010011100100001011000" , -- ADDR 1041
			"00000000000010001000011110101001" , -- ADDR 1042
			"00000000000011000101101000000011" , -- ADDR 1043
			"00000000000001101000100111100011" , -- ADDR 1044
			"00000000000001010100000101100100" , -- ADDR 1045
			"00000000000001110010101001000110" , -- ADDR 1046
			"00000000000010100110110001101110" , -- ADDR 1047
			"00000000000010100000001101011100" , -- ADDR 1048
			"00000000000001010010010101001111" , -- ADDR 1049
			"00000000000001111101011110001011" , -- ADDR 1050
			"00000000000000111111011000011111" , -- ADDR 1051
			"00000000000001101100101100101001" , -- ADDR 1052
			"00000000000001111000001101101000" , -- ADDR 1053
			"00000000000100001011011111111001" , -- ADDR 1054
			"00000000000001100010001001001011" , -- ADDR 1055
			"00000000000001100101100000001000" , -- ADDR 1056
			"00000000000001101001001010000110" , -- ADDR 1057
			"00000000000001101100010111000111" , -- ADDR 1058
			"00000000000001110110001101101000" , -- ADDR 1059
			"00000000000001110000000010111011" , -- ADDR 1060
			"00000000000001110101010100001001" , -- ADDR 1061
			"00000000000011000011101101100111" , -- ADDR 1062
			"00000000000010001011010100001100" , -- ADDR 1063
			"00000000000010111100001000101000" , -- ADDR 1064
			"00000000000001001110101110111010" , -- ADDR 1065
			"00000000000010011101001000100111" , -- ADDR 1066
			"00000000000001010101001111111010" , -- ADDR 1067
			"00000000000001111111101000110101" , -- ADDR 1068
			"00000000000001110000111000110001" , -- ADDR 1069
			"00000000000001101101011110000010" , -- ADDR 1070
			"00000000000000101110101110010001" , -- ADDR 1071
			"00000000000011010100110000011010" , -- ADDR 1072
			"00000000000100001000001001100010" , -- ADDR 1073
			"00000000000001001010100000001100" , -- ADDR 1074
			"00000000000001101101000010000110" , -- ADDR 1075
			"00000000000100011110010110100110" , -- ADDR 1076
			"00000000000001101011010000010110" , -- ADDR 1077
			"00000000000001101011101101101000" , -- ADDR 1078
			"00000000000001101110100110011010" , -- ADDR 1079
			"00000000000001111100010010111101" , -- ADDR 1080
			"00000000000010000110101010100101" , -- ADDR 1081
			"00000000000001111000101011010100" , -- ADDR 1082
			"00000000000010000001110000110011" , -- ADDR 1083
			"00000000000010101110000100001001" , -- ADDR 1084
			"00000000000001001100111100010111" , -- ADDR 1085
			"00000000000011000111000111000000" , -- ADDR 1086
			"00000000000001011101011110100100" , -- ADDR 1087
			"00000000000010001110011010001110" , -- ADDR 1088
			"00000000000001110101011111111010" , -- ADDR 1089
			"00000000000010111110111101110000" , -- ADDR 1090
			"00000000000010000111000011010101" , -- ADDR 1091
			"00000000000001100111001100001110" , -- ADDR 1092
			"00000000000000110100100011000000" , -- ADDR 1093
			"00000000000011111110111100111010" , -- ADDR 1094
			"00000000000101000100101101011001" , -- ADDR 1095
			"00000000000000101110011001110010" , -- ADDR 1096
			"00000000000011100111011110010101" , -- ADDR 1097
			"00000000000001000100101000011010" , -- ADDR 1098
			"00000000000001000001011011100010" , -- ADDR 1099
			"00000000000001000010000100110111" , -- ADDR 1100
			"00000000000001010110011111110111" , -- ADDR 1101
			"00000000000001011110001001110001" , -- ADDR 1102
			"00000000000001001011110011010011" , -- ADDR 1103
			"00000000000001010110001011111111" , -- ADDR 1104
			"00000000000001100011110010001110" , -- ADDR 1105
			"00000000000001101011001010000111" , -- ADDR 1106
			"00000000000010001110011010001110" , -- ADDR 1107
			"00000000000001000101101010100111" , -- ADDR 1108
			"00000000000001000111100001011111" , -- ADDR 1109
			"00000000000001100101100010111101" , -- ADDR 1110
			"00000000000011011010101110000111" , -- ADDR 1111
			"00000000000001100100111111101001" , -- ADDR 1112
			"00000000000000110000010010101000" , -- ADDR 1113
			"00000000000000111111111101111011" , -- ADDR 1114
			"00000000000011100100011010010111" , -- ADDR 1115
			"00000000000101001011000010001001" , -- ADDR 1116
			"00000000000010111001001110111100" , -- ADDR 1117
			"00000000000000100100111001111010" , -- ADDR 1118
			"00000000000000011111110101010000" , -- ADDR 1119
			"00000000000000011110000001101000" , -- ADDR 1120
			"00000000000000110001011101110000" , -- ADDR 1121
			"00000000000000110101111011101011" , -- ADDR 1122
			"00000000000000100100001001100111" , -- ADDR 1123
			"00000000000000101101010100000111" , -- ADDR 1124
			"00000000000001001100000011000000" , -- ADDR 1125
			"00000000000010011001010101000001" , -- ADDR 1126
			"00000000000001100000001000000100" , -- ADDR 1127
			"00000000000000110010100010011010" , -- ADDR 1128
			"00000000000000100100111100011111" , -- ADDR 1129
			"00000000000001001100001101000010" , -- ADDR 1130
			"00000000000011001110010011001000" , -- ADDR 1131
			"00000000000000111111101100000000" , -- ADDR 1132
			"00000000000000001100001101010000" , -- ADDR 1133
			"00000000000001001010100111110111" , -- ADDR 1134
			"00000000000010111011010101110101" , -- ADDR 1135
			"00000000000100101110010101111100" , -- ADDR 1136
			"00000000000010110011001110010010" , -- ADDR 1137
			"00000000000010110010101001100000" , -- ADDR 1138
			"00000000000010101111110101100010" , -- ADDR 1139
			"00000000000010100011001101011010" , -- ADDR 1140
			"00000000000010011000101101011100" , -- ADDR 1141
			"00000000000010100101101011011100" , -- ADDR 1142
			"00000000000010011100101111101100" , -- ADDR 1143
			"00000000000010101011111000000110" , -- ADDR 1144
			"00000000000101010010100011101100" , -- ADDR 1145
			"00000000000001011001000111001000" , -- ADDR 1146
			"00000000000011000011000001011100" , -- ADDR 1147
			"00000000000010100111111010101010" , -- ADDR 1148
			"00000000000010110110011000000011" , -- ADDR 1149
			"00000000000100001011011000001111" , -- ADDR 1150
			"00000000000010011011010110011110" , -- ADDR 1151
			"00000000000010111010011100111100" , -- ADDR 1152
			"00000000000011101101101101100010" , -- ADDR 1153
			"00000000000001110011111000111100" , -- ADDR 1154
			"00000000000100001001110011010110" , -- ADDR 1155
			"00000000000000000101001011011101" , -- ADDR 1156
			"00000000000000001000001100000101" , -- ADDR 1157
			"00000000000000010010100101111110" , -- ADDR 1158
			"00000000000000011100000110100101" , -- ADDR 1159
			"00000000000000001110010010011011" , -- ADDR 1160
			"00000000000000010110100000100011" , -- ADDR 1161
			"00000000000001101011110100010000" , -- ADDR 1162
			"00000000000010100111000110000000" , -- ADDR 1163
			"00000000000001011101010110111010" , -- ADDR 1164
			"00000000000000010011100010000000" , -- ADDR 1165
			"00000000000001000011011010100110" , -- ADDR 1166
			"00000000000000100111010011110100" , -- ADDR 1167
			"00000000000010101010001110001011" , -- ADDR 1168
			"00000000000000100000100100101001" , -- ADDR 1169
			"00000000000000011001101010011111" , -- ADDR 1170
			"00000000000000111011100000111100" , -- ADDR 1171
			"00000000000010100000001101011100" , -- ADDR 1172
			"00000000000100001010110000001111" , -- ADDR 1173
			"00000000000000000011101010011000" , -- ADDR 1174
			"00000000000000010101000100101001" , -- ADDR 1175
			"00000000000000011101011111111110" , -- ADDR 1176
			"00000000000000001100111110011111" , -- ADDR 1177
			"00000000000000010110101101001101" , -- ADDR 1178
			"00000000000001100110110011101100" , -- ADDR 1179
			"00000000000010100101101001001001" , -- ADDR 1180
			"00000000000001011011111010010000" , -- ADDR 1181
			"00000000000000010111011110110001" , -- ADDR 1182
			"00000000000000111110011000110011" , -- ADDR 1183
			"00000000000000101100011011110011" , -- ADDR 1184
			"00000000000010101111011001010010" , -- ADDR 1185
			"00000000000000100011100101101110" , -- ADDR 1186
			"00000000000000010100110111000000" , -- ADDR 1187
			"00000000000000111101011011111101" , -- ADDR 1188
			"00000000000010100011000010000000" , -- ADDR 1189
			"00000000000100001111010111110110" , -- ADDR 1190
			"00000000000000010100110000001000" , -- ADDR 1191
			"00000000000000011100001011101010" , -- ADDR 1192
			"00000000000000001010100000000100" , -- ADDR 1193
			"00000000000000010100110000001000" , -- ADDR 1194
			"00000000000001100011101001100111" , -- ADDR 1195
			"00000000000010100111011110110011" , -- ADDR 1196
			"00000000000001011000110001001001" , -- ADDR 1197
			"00000000000000011011000110101010" , -- ADDR 1198
			"00000000000000111011010000111001" , -- ADDR 1199
			"00000000000000101110101111010010" , -- ADDR 1200
			"00000000000010110010000111010011" , -- ADDR 1201
			"00000000000000100011011001101000" , -- ADDR 1202
			"00000000000000010011110111110010" , -- ADDR 1203
			"00000000000001000000110111101011" , -- ADDR 1204
			"00000000000010100010010110111011" , -- ADDR 1205
			"00000000000100010000100011000100" , -- ADDR 1206
			"00000000000000001010100000000100" , -- ADDR 1207
			"00000000000000001101101001011110" , -- ADDR 1208
			"00000000000000001010000100001111" , -- ADDR 1209
			"00000000000001101111110000001011" , -- ADDR 1210
			"00000000000010111001101000011001" , -- ADDR 1211
			"00000000000001001111111010000100" , -- ADDR 1212
			"00000000000000011111110101010000" , -- ADDR 1213
			"00000000000001001000100001101101" , -- ADDR 1214
			"00000000000000100001110110011110" , -- ADDR 1215
			"00000000000010100101000011000100" , -- ADDR 1216
			"00000000000000001110101001100000" , -- ADDR 1217
			"00000000000000101000011100110000" , -- ADDR 1218
			"00000000000001001010100000001100" , -- ADDR 1219
			"00000000000010001101111101101101" , -- ADDR 1220
			"00000000000011111101000001110000" , -- ADDR 1221
			"00000000000000010010011110010000" , -- ADDR 1222
			"00000000000000001000101000011011" , -- ADDR 1223
			"00000000000001101101101000000011" , -- ADDR 1224
			"00000000000011000011000010101010" , -- ADDR 1225
			"00000000000001000101111011000000" , -- ADDR 1226
			"00000000000000101010010100100101" , -- ADDR 1227
			"00000000000001000111110011011101" , -- ADDR 1228
			"00000000000000100111111111000111" , -- ADDR 1229
			"00000000000010101000100111101110" , -- ADDR 1230
			"00000000000000001100000101011001" , -- ADDR 1231
			"00000000000000101110101001001010" , -- ADDR 1232
			"00000000000001010101000000001110" , -- ADDR 1233
			"00000000000010000110011110111000" , -- ADDR 1234
			"00000000000011111010100001111010" , -- ADDR 1235
			"00000000000000001010011011100000" , -- ADDR 1236
			"00000000000001100011010111011001" , -- ADDR 1237
			"00000000000010110001111100100101" , -- ADDR 1238
			"00000000000001001111001101000111" , -- ADDR 1239
			"00000000000000100001010100011001" , -- ADDR 1240
			"00000000000000111011100111010110" , -- ADDR 1241
			"00000000000000101101011010011011" , -- ADDR 1242
			"00000000000010110001010011001111" , -- ADDR 1243
			"00000000000000011011100010100101" , -- ADDR 1244
			"00000000000000011100001011101010" , -- ADDR 1245
			"00000000000001001001101111111100" , -- ADDR 1246
			"00000000000010011000111101000010" , -- ADDR 1247
			"00000000000100001010100110110000" , -- ADDR 1248
			"00000000000001100110110011101100" , -- ADDR 1249
			"00000000000010111100001101101101" , -- ADDR 1250
			"00000000000001000111101001011111" , -- ADDR 1251
			"00000000000000100111011100010011" , -- ADDR 1252
			"00000000000001000000001111110010" , -- ADDR 1253
			"00000000000000101011110000100010" , -- ADDR 1254
			"00000000000010101110011010000010" , -- ADDR 1255
			"00000000000000010011101011101111" , -- ADDR 1256
			"00000000000000100110010101001011" , -- ADDR 1257
			"00000000000001010001011101010110" , -- ADDR 1258
			"00000000000010001110110001111101" , -- ADDR 1259
			"00000000000100000010111000100101" , -- ADDR 1260
			"00000000000011000010011101001100" , -- ADDR 1261
			"00000000000001100010001001001011" , -- ADDR 1262
			"00000000000001111101000001001111" , -- ADDR 1263
			"00000000000000101000011011100101" , -- ADDR 1264
			"00000000000010010000110001101001" , -- ADDR 1265
			"00000000000100010100101001100111" , -- ADDR 1266
			"00000000000001111001101101011011" , -- ADDR 1267
			"00000000000001010111101110101100" , -- ADDR 1268
			"00000000000010010101011000101010" , -- ADDR 1269
			"00000000000011011010110101100010" , -- ADDR 1270
			"00000000000101100010110000011011" , -- ADDR 1271
			"00000000000011111001011101000011" , -- ADDR 1272
			"00000000000010011110111001110001" , -- ADDR 1273
			"00000000000010101111111111010010" , -- ADDR 1274
			"00000000000010111011101010011100" , -- ADDR 1275
			"00000000000100001010101110111111" , -- ADDR 1276
			"00000000000011000110101111111111" , -- ADDR 1277
			"00000000000010011001000111010100" , -- ADDR 1278
			"00000000000001111100011111001110" , -- ADDR 1279
			"00000000000101000100011101101011" , -- ADDR 1280
			"00000000000110010001101000001100" , -- ADDR 1281
			"00000000000001101111000101011000" , -- ADDR 1282
			"00000000000001010010001110010010" , -- ADDR 1283
			"00000000000001101010110001001001" , -- ADDR 1284
			"00000000000011011100110100001101" , -- ADDR 1285
			"00000000000001001100011110100001" , -- ADDR 1286
			"00000000000001100001101000100010" , -- ADDR 1287
			"00000000000010011000110110110011" , -- ADDR 1288
			"00000000000001111011000110101000" , -- ADDR 1289
			"00000000000100001011110111110001" , -- ADDR 1290
			"00000000000001010100101010010011" , -- ADDR 1291
			"00000000000000011111111100101111" , -- ADDR 1292
			"00000000000010011100010110011010" , -- ADDR 1293
			"00000000000000101001100100110110" , -- ADDR 1294
			"00000000000000100110010101001011" , -- ADDR 1295
			"00000000000000101010101110011000" , -- ADDR 1296
			"00000000000010100101100111111111" , -- ADDR 1297
			"00000000000100000101011011010110" , -- ADDR 1298
			"00000000000001101000110111111100" , -- ADDR 1299
			"00000000000011101100110010110110" , -- ADDR 1300
			"00000000000001010011101111011001" , -- ADDR 1301
			"00000000000000101111111101110101" , -- ADDR 1302
			"00000000000001101111100000110011" , -- ADDR 1303
			"00000000000011000000111001111110" , -- ADDR 1304
			"00000000000101000001000010010010" , -- ADDR 1305
			"00000000000010000011111011010010" , -- ADDR 1306
			"00000000000000011110100001001000" , -- ADDR 1307
			"00000000000001000000101100101000" , -- ADDR 1308
			"00000000000001000000111111000001" , -- ADDR 1309
			"00000000000010001001100111000001" , -- ADDR 1310
			"00000000000011100101110000111100" , -- ADDR 1311
			"00000000000010011100110100110111" , -- ADDR 1312
			"00000000000011000010001101101111" , -- ADDR 1313
			"00000000000010011101110001110010" , -- ADDR 1314
			"00000000000010100110011001000110" , -- ADDR 1315
			"00000000000010010001111011110010" , -- ADDR 1316
			"00000000000000110111000011011011" , -- ADDR 1317
			"00000000000001010011110001000111" , -- ADDR 1318
			"00000000000001111111101000110101" , -- ADDR 1319
			"00000000000011101111010111111000" , -- ADDR 1320
			"00000000000001000000101111100101" , -- ADDR 1321
			"00000000000010110101000110001100" , -- ADDR 1322
			"00000000000100100100001101111011" , -- ADDR 1323
			"00000000000011001010100010101000" , -- ADDR 1324
			"00000000000100011000111100101001" , -- ADDR 1325
			"00000000000010011000100010110100" , -- ADDR 1326
			"00000000000000000000000000000000" , -- ADDR 1327
			"00000000000000000000000000000000" , -- ADDR 1328
			"00000000000000000000000000000000" , -- ADDR 1329
			"00000000000000000000000000000000" , -- ADDR 1330
			"00000000000000000000000000000000" , -- ADDR 1331
			"00000000000000000000000000000000" , -- ADDR 1332
			"00000000000000000000000000000000" , -- ADDR 1333
			"00000000000000000000000000000000" , -- ADDR 1334
			"00000000000000000000000000000000" , -- ADDR 1335
			"00000000000000000000000000000000" , -- ADDR 1336
			"00000000000000000000000000000000" , -- ADDR 1337
			"00000000000000000000000000000000" , -- ADDR 1338
			"00000000000000000000000000000000" , -- ADDR 1339
			"00000000000000000000000000000000" , -- ADDR 1340
			"00000000000000000000000000000000" , -- ADDR 1341
			"00000000000000000000000000000000" , -- ADDR 1342
			"00000000000000000000000000000000" , -- ADDR 1343
			"00000000000000000000000000000000" , -- ADDR 1344
			"00000000000000000000000000000000" , -- ADDR 1345
			"00000000000000000000000000000000" , -- ADDR 1346
			"00000000000000000000000000000000" , -- ADDR 1347
			"00000000000000000000000000000000" , -- ADDR 1348
			"00000000000000000000000000000000" , -- ADDR 1349
			"00000000000000000000000000000000" , -- ADDR 1350
			"00000000000000000000000000000000" , -- ADDR 1351
			"00000000000000000000000000000000" , -- ADDR 1352
			"00000000000000000000000000000000" , -- ADDR 1353
			"00000000000000000000000000000000" , -- ADDR 1354
			"00000000000000000000000000000000" , -- ADDR 1355
			"00000000000000000000000000000000" , -- ADDR 1356
			"00000000000000000000000000000000" , -- ADDR 1357
			"00000000000000000000000000000000" , -- ADDR 1358
			"00000000000000000000000000000000" , -- ADDR 1359
			"00000000000000000000000000000000" , -- ADDR 1360
			"00000000000000000000000000000000" , -- ADDR 1361
			"00000000000000000000000000000000" , -- ADDR 1362
			"00000000000000000000000000000000" , -- ADDR 1363
			"00000000000000000000000000000000" , -- ADDR 1364
			"00000000000000000000000000000000" , -- ADDR 1365
			"00000000000000000000000000000000" , -- ADDR 1366
			"00000000000000000000000000000000" , -- ADDR 1367
			"00000000000000000000000000000000" , -- ADDR 1368
			"00000000000000000000000000000000" , -- ADDR 1369
			"00000000000000000000000000000000" , -- ADDR 1370
			"00000000000000000000000000000000" , -- ADDR 1371
			"00000000000000000000000000000000" , -- ADDR 1372
			"00000000000000000000000000000000" , -- ADDR 1373
			"00000000000000000000000000000000" , -- ADDR 1374
			"00000000000000000000000000000000" , -- ADDR 1375
			"00000000000000000000000000000000" , -- ADDR 1376
			"00000000000000000000000000000000" , -- ADDR 1377
			"00000000000000000000000000000000" , -- ADDR 1378
			"00000000000000000000000000000000" , -- ADDR 1379
			"00000000000000000000000000000000" , -- ADDR 1380
			"00000000000000000000000000000000" , -- ADDR 1381
			"00000000000000000000000000000000" , -- ADDR 1382
			"00000000000000000000000000000000" , -- ADDR 1383
			"00000000000000000000000000000000" , -- ADDR 1384
			"00000000000000000000000000000000" , -- ADDR 1385
			"00000000000000000000000000000000" , -- ADDR 1386
			"00000000000000000000000000000000" , -- ADDR 1387
			"00000000000000000000000000000000" , -- ADDR 1388
			"00000000000000000000000000000000" , -- ADDR 1389
			"00000000000000000000000000000000" , -- ADDR 1390
			"00000000000000000000000000000000" , -- ADDR 1391
			"00000000000000000000000000000000" , -- ADDR 1392
			"00000000000000000000000000000000" , -- ADDR 1393
			"00000000000000000000000000000000" , -- ADDR 1394
			"00000000000000000000000000000000" , -- ADDR 1395
			"00000000000000000000000000000000" , -- ADDR 1396
			"00000000000000000000000000000000" , -- ADDR 1397
			"00000000000000000000000000000000" , -- ADDR 1398
			"00000000000000000000000000000000" , -- ADDR 1399
			"00000000000000000000000000000000" , -- ADDR 1400
			"00000000000000000000000000000000" , -- ADDR 1401
			"00000000000000000000000000000000" , -- ADDR 1402
			"00000000000000000000000000000000" , -- ADDR 1403
			"00000000000000000000000000000000" , -- ADDR 1404
			"00000000000000000000000000000000" , -- ADDR 1405
			"00000000000000000000000000000000" , -- ADDR 1406
			"00000000000000000000000000000000" , -- ADDR 1407
			"00000000000000000000000000000000" , -- ADDR 1408
			"00000000000000000000000000000000" , -- ADDR 1409
			"00000000000000000000000000000000" , -- ADDR 1410
			"00000000000000000000000000000000" , -- ADDR 1411
			"00000000000000000000000000000000" , -- ADDR 1412
			"00000000000000000000000000000000" , -- ADDR 1413
			"00000000000000000000000000000000" , -- ADDR 1414
			"00000000000000000000000000000000" , -- ADDR 1415
			"00000000000000000000000000000000" , -- ADDR 1416
			"00000000000000000000000000000000" , -- ADDR 1417
			"00000000000000000000000000000000" , -- ADDR 1418
			"00000000000000000000000000000000" , -- ADDR 1419
			"00000000000000000000000000000000" , -- ADDR 1420
			"00000000000000000000000000000000" , -- ADDR 1421
			"00000000000000000000000000000000" , -- ADDR 1422
			"00000000000000000000000000000000" , -- ADDR 1423
			"00000000000000000000000000000000" , -- ADDR 1424
			"00000000000000000000000000000000" , -- ADDR 1425
			"00000000000000000000000000000000" , -- ADDR 1426
			"00000000000000000000000000000000" , -- ADDR 1427
			"00000000000000000000000000000000" , -- ADDR 1428
			"00000000000000000000000000000000" , -- ADDR 1429
			"00000000000000000000000000000000" , -- ADDR 1430
			"00000000000000000000000000000000" , -- ADDR 1431
			"00000000000000000000000000000000" , -- ADDR 1432
			"00000000000000000000000000000000" , -- ADDR 1433
			"00000000000000000000000000000000" , -- ADDR 1434
			"00000000000000000000000000000000" , -- ADDR 1435
			"00000000000000000000000000000000" , -- ADDR 1436
			"00000000000000000000000000000000" , -- ADDR 1437
			"00000000000000000000000000000000" , -- ADDR 1438
			"00000000000000000000000000000000" , -- ADDR 1439
			"00000000000000000000000000000000" , -- ADDR 1440
			"00000000000000000000000000000000" , -- ADDR 1441
			"00000000000000000000000000000000" , -- ADDR 1442
			"00000000000000000000000000000000" , -- ADDR 1443
			"00000000000000000000000000000000" , -- ADDR 1444
			"00000000000000000000000000000000" , -- ADDR 1445
			"00000000000000000000000000000000" , -- ADDR 1446
			"00000000000000000000000000000000" , -- ADDR 1447
			"00000000000000000000000000000000" , -- ADDR 1448
			"00000000000000000000000000000000" , -- ADDR 1449
			"00000000000000000000000000000000" , -- ADDR 1450
			"00000000000000000000000000000000" , -- ADDR 1451
			"00000000000000000000000000000000" , -- ADDR 1452
			"00000000000000000000000000000000" , -- ADDR 1453
			"00000000000000000000000000000000" , -- ADDR 1454
			"00000000000000000000000000000000" , -- ADDR 1455
			"00000000000000000000000000000000" , -- ADDR 1456
			"00000000000000000000000000000000" , -- ADDR 1457
			"00000000000000000000000000000000" , -- ADDR 1458
			"00000000000000000000000000000000" , -- ADDR 1459
			"00000000000000000000000000000000" , -- ADDR 1460
			"00000000000000000000000000000000" , -- ADDR 1461
			"00000000000000000000000000000000" , -- ADDR 1462
			"00000000000000000000000000000000" , -- ADDR 1463
			"00000000000000000000000000000000" , -- ADDR 1464
			"00000000000000000000000000000000" , -- ADDR 1465
			"00000000000000000000000000000000" , -- ADDR 1466
			"00000000000000000000000000000000" , -- ADDR 1467
			"00000000000000000000000000000000" , -- ADDR 1468
			"00000000000000000000000000000000" , -- ADDR 1469
			"00000000000000000000000000000000" , -- ADDR 1470
			"00000000000000000000000000000000" , -- ADDR 1471
			"00000000000000000000000000000000" , -- ADDR 1472
			"00000000000000000000000000000000" , -- ADDR 1473
			"00000000000000000000000000000000" , -- ADDR 1474
			"00000000000000000000000000000000" , -- ADDR 1475
			"00000000000000000000000000000000" , -- ADDR 1476
			"00000000000000000000000000000000" , -- ADDR 1477
			"00000000000000000000000000000000" , -- ADDR 1478
			"00000000000000000000000000000000" , -- ADDR 1479
			"00000000000000000000000000000000" , -- ADDR 1480
			"00000000000000000000000000000000" , -- ADDR 1481
			"00000000000000000000000000000000" , -- ADDR 1482
			"00000000000000000000000000000000" , -- ADDR 1483
			"00000000000000000000000000000000" , -- ADDR 1484
			"00000000000000000000000000000000" , -- ADDR 1485
			"00000000000000000000000000000000" , -- ADDR 1486
			"00000000000000000000000000000000" , -- ADDR 1487
			"00000000000000000000000000000000" , -- ADDR 1488
			"00000000000000000000000000000000" , -- ADDR 1489
			"00000000000000000000000000000000" , -- ADDR 1490
			"00000000000000000000000000000000" , -- ADDR 1491
			"00000000000000000000000000000000" , -- ADDR 1492
			"00000000000000000000000000000000" , -- ADDR 1493
			"00000000000000000000000000000000" , -- ADDR 1494
			"00000000000000000000000000000000" , -- ADDR 1495
			"00000000000000000000000000000000" , -- ADDR 1496
			"00000000000000000000000000000000" , -- ADDR 1497
			"00000000000000000000000000000000" , -- ADDR 1498
			"00000000000000000000000000000000" , -- ADDR 1499
			"00000000000000000000000000000000" , -- ADDR 1500
			"00000000000000000000000000000000" , -- ADDR 1501
			"00000000000000000000000000000000" , -- ADDR 1502
			"00000000000000000000000000000000" , -- ADDR 1503
			"00000000000000000000000000000000" , -- ADDR 1504
			"00000000000000000000000000000000" , -- ADDR 1505
			"00000000000000000000000000000000" , -- ADDR 1506
			"00000000000000000000000000000000" , -- ADDR 1507
			"00000000000000000000000000000000" , -- ADDR 1508
			"00000000000000000000000000000000" , -- ADDR 1509
			"00000000000000000000000000000000" , -- ADDR 1510
			"00000000000000000000000000000000" , -- ADDR 1511
			"00000000000000000000000000000000" , -- ADDR 1512
			"00000000000000000000000000000000" , -- ADDR 1513
			"00000000000000000000000000000000" , -- ADDR 1514
			"00000000000000000000000000000000" , -- ADDR 1515
			"00000000000000000000000000000000" , -- ADDR 1516
			"00000000000000000000000000000000" , -- ADDR 1517
			"00000000000000000000000000000000" , -- ADDR 1518
			"00000000000000000000000000000000" , -- ADDR 1519
			"00000000000000000000000000000000" , -- ADDR 1520
			"00000000000000000000000000000000" , -- ADDR 1521
			"00000000000000000000000000000000" , -- ADDR 1522
			"00000000000000000000000000000000" , -- ADDR 1523
			"00000000000000000000000000000000" , -- ADDR 1524
			"00000000000000000000000000000000" , -- ADDR 1525
			"00000000000000000000000000000000" , -- ADDR 1526
			"00000000000000000000000000000000" , -- ADDR 1527
			"00000000000000000000000000000000" , -- ADDR 1528
			"00000000000000000000000000000000" , -- ADDR 1529
			"00000000000000000000000000000000" , -- ADDR 1530
			"00000000000000000000000000000000" , -- ADDR 1531
			"00000000000000000000000000000000" , -- ADDR 1532
			"00000000000000000000000000000000" , -- ADDR 1533
			"00000000000000000000000000000000" , -- ADDR 1534
			"00000000000000000000000000000000" , -- ADDR 1535
			"00000000000000000000000000000000" , -- ADDR 1536
			"00000000000000000000000000000000" , -- ADDR 1537
			"00000000000000000000000000000000" , -- ADDR 1538
			"00000000000000000000000000000000" , -- ADDR 1539
			"00000000000000000000000000000000" , -- ADDR 1540
			"00000000000000000000000000000000" , -- ADDR 1541
			"00000000000000000000000000000000" , -- ADDR 1542
			"00000000000000000000000000000000" , -- ADDR 1543
			"00000000000000000000000000000000" , -- ADDR 1544
			"00000000000000000000000000000000" , -- ADDR 1545
			"00000000000000000000000000000000" , -- ADDR 1546
			"00000000000000000000000000000000" , -- ADDR 1547
			"00000000000000000000000000000000" , -- ADDR 1548
			"00000000000000000000000000000000" , -- ADDR 1549
			"00000000000000000000000000000000" , -- ADDR 1550
			"00000000000000000000000000000000" , -- ADDR 1551
			"00000000000000000000000000000000" , -- ADDR 1552
			"00000000000000000000000000000000" , -- ADDR 1553
			"00000000000000000000000000000000" , -- ADDR 1554
			"00000000000000000000000000000000" , -- ADDR 1555
			"00000000000000000000000000000000" , -- ADDR 1556
			"00000000000000000000000000000000" , -- ADDR 1557
			"00000000000000000000000000000000" , -- ADDR 1558
			"00000000000000000000000000000000" , -- ADDR 1559
			"00000000000000000000000000000000" , -- ADDR 1560
			"00000000000000000000000000000000" , -- ADDR 1561
			"00000000000000000000000000000000" , -- ADDR 1562
			"00000000000000000000000000000000" , -- ADDR 1563
			"00000000000000000000000000000000" , -- ADDR 1564
			"00000000000000000000000000000000" , -- ADDR 1565
			"00000000000000000000000000000000" , -- ADDR 1566
			"00000000000000000000000000000000" , -- ADDR 1567
			"00000000000000000000000000000000" , -- ADDR 1568
			"00000000000000000000000000000000" , -- ADDR 1569
			"00000000000000000000000000000000" , -- ADDR 1570
			"00000000000000000000000000000000" , -- ADDR 1571
			"00000000000000000000000000000000" , -- ADDR 1572
			"00000000000000000000000000000000" , -- ADDR 1573
			"00000000000000000000000000000000" , -- ADDR 1574
			"00000000000000000000000000000000" , -- ADDR 1575
			"00000000000000000000000000000000" , -- ADDR 1576
			"00000000000000000000000000000000" , -- ADDR 1577
			"00000000000000000000000000000000" , -- ADDR 1578
			"00000000000000000000000000000000" , -- ADDR 1579
			"00000000000000000000000000000000" , -- ADDR 1580
			"00000000000000000000000000000000" , -- ADDR 1581
			"00000000000000000000000000000000" , -- ADDR 1582
			"00000000000000000000000000000000" , -- ADDR 1583
			"00000000000000000000000000000000" , -- ADDR 1584
			"00000000000000000000000000000000" , -- ADDR 1585
			"00000000000000000000000000000000" , -- ADDR 1586
			"00000000000000000000000000000000" , -- ADDR 1587
			"00000000000000000000000000000000" , -- ADDR 1588
			"00000000000000000000000000000000" , -- ADDR 1589
			"00000000000000000000000000000000" , -- ADDR 1590
			"00000000000000000000000000000000" , -- ADDR 1591
			"00000000000000000000000000000000" , -- ADDR 1592
			"00000000000000000000000000000000" , -- ADDR 1593
			"00000000000000000000000000000000" , -- ADDR 1594
			"00000000000000000000000000000000" , -- ADDR 1595
			"00000000000000000000000000000000" , -- ADDR 1596
			"00000000000000000000000000000000" , -- ADDR 1597
			"00000000000000000000000000000000" , -- ADDR 1598
			"00000000000000000000000000000000" , -- ADDR 1599
			"00000000000000000000000000000000" , -- ADDR 1600
			"00000000000000000000000000000000" , -- ADDR 1601
			"00000000000000000000000000000000" , -- ADDR 1602
			"00000000000000000000000000000000" , -- ADDR 1603
			"00000000000000000000000000000000" , -- ADDR 1604
			"00000000000000000000000000000000" , -- ADDR 1605
			"00000000000000000000000000000000" , -- ADDR 1606
			"00000000000000000000000000000000" , -- ADDR 1607
			"00000000000000000000000000000000" , -- ADDR 1608
			"00000000000000000000000000000000" , -- ADDR 1609
			"00000000000000000000000000000000" , -- ADDR 1610
			"00000000000000000000000000000000" , -- ADDR 1611
			"00000000000000000000000000000000" , -- ADDR 1612
			"00000000000000000000000000000000" , -- ADDR 1613
			"00000000000000000000000000000000" , -- ADDR 1614
			"00000000000000000000000000000000" , -- ADDR 1615
			"00000000000000000000000000000000" , -- ADDR 1616
			"00000000000000000000000000000000" , -- ADDR 1617
			"00000000000000000000000000000000" , -- ADDR 1618
			"00000000000000000000000000000000" , -- ADDR 1619
			"00000000000000000000000000000000" , -- ADDR 1620
			"00000000000000000000000000000000" , -- ADDR 1621
			"00000000000000000000000000000000" , -- ADDR 1622
			"00000000000000000000000000000000" , -- ADDR 1623
			"00000000000000000000000000000000" , -- ADDR 1624
			"00000000000000000000000000000000" , -- ADDR 1625
			"00000000000000000000000000000000" , -- ADDR 1626
			"00000000000000000000000000000000" , -- ADDR 1627
			"00000000000000000000000000000000" , -- ADDR 1628
			"00000000000000000000000000000000" , -- ADDR 1629
			"00000000000000000000000000000000" , -- ADDR 1630
			"00000000000000000000000000000000" , -- ADDR 1631
			"00000000000000000000000000000000" , -- ADDR 1632
			"00000000000000000000000000000000" , -- ADDR 1633
			"00000000000000000000000000000000" , -- ADDR 1634
			"00000000000000000000000000000000" , -- ADDR 1635
			"00000000000000000000000000000000" , -- ADDR 1636
			"00000000000000000000000000000000" , -- ADDR 1637
			"00000000000000000000000000000000" , -- ADDR 1638
			"00000000000000000000000000000000" , -- ADDR 1639
			"00000000000000000000000000000000" , -- ADDR 1640
			"00000000000000000000000000000000" , -- ADDR 1641
			"00000000000000000000000000000000" , -- ADDR 1642
			"00000000000000000000000000000000" , -- ADDR 1643
			"00000000000000000000000000000000" , -- ADDR 1644
			"00000000000000000000000000000000" , -- ADDR 1645
			"00000000000000000000000000000000" , -- ADDR 1646
			"00000000000000000000000000000000" , -- ADDR 1647
			"00000000000000000000000000000000" , -- ADDR 1648
			"00000000000000000000000000000000" , -- ADDR 1649
			"00000000000000000000000000000000" , -- ADDR 1650
			"00000000000000000000000000000000" , -- ADDR 1651
			"00000000000000000000000000000000" , -- ADDR 1652
			"00000000000000000000000000000000" , -- ADDR 1653
			"00000000000000000000000000000000" , -- ADDR 1654
			"00000000000000000000000000000000" , -- ADDR 1655
			"00000000000000000000000000000000" , -- ADDR 1656
			"00000000000000000000000000000000" , -- ADDR 1657
			"00000000000000000000000000000000" , -- ADDR 1658
			"00000000000000000000000000000000" , -- ADDR 1659
			"00000000000000000000000000000000" , -- ADDR 1660
			"00000000000000000000000000000000" , -- ADDR 1661
			"00000000000000000000000000000000" , -- ADDR 1662
			"00000000000000000000000000000000" , -- ADDR 1663
			"00000000000000000000000000000000" , -- ADDR 1664
			"00000000000000000000000000000000" , -- ADDR 1665
			"00000000000000000000000000000000" , -- ADDR 1666
			"00000000000000000000000000000000" , -- ADDR 1667
			"00000000000000000000000000000000" , -- ADDR 1668
			"00000000000000000000000000000000" , -- ADDR 1669
			"00000000000000000000000000000000" , -- ADDR 1670
			"00000000000000000000000000000000" , -- ADDR 1671
			"00000000000000000000000000000000" , -- ADDR 1672
			"00000000000000000000000000000000" , -- ADDR 1673
			"00000000000000000000000000000000" , -- ADDR 1674
			"00000000000000000000000000000000" , -- ADDR 1675
			"00000000000000000000000000000000" , -- ADDR 1676
			"00000000000000000000000000000000" , -- ADDR 1677
			"00000000000000000000000000000000" , -- ADDR 1678
			"00000000000000000000000000000000" , -- ADDR 1679
			"00000000000000000000000000000000" , -- ADDR 1680
			"00000000000000000000000000000000" , -- ADDR 1681
			"00000000000000000000000000000000" , -- ADDR 1682
			"00000000000000000000000000000000" , -- ADDR 1683
			"00000000000000000000000000000000" , -- ADDR 1684
			"00000000000000000000000000000000" , -- ADDR 1685
			"00000000000000000000000000000000" , -- ADDR 1686
			"00000000000000000000000000000000" , -- ADDR 1687
			"00000000000000000000000000000000" , -- ADDR 1688
			"00000000000000000000000000000000" , -- ADDR 1689
			"00000000000000000000000000000000" , -- ADDR 1690
			"00000000000000000000000000000000" , -- ADDR 1691
			"00000000000000000000000000000000" , -- ADDR 1692
			"00000000000000000000000000000000" , -- ADDR 1693
			"00000000000000000000000000000000" , -- ADDR 1694
			"00000000000000000000000000000000" , -- ADDR 1695
			"00000000000000000000000000000000" , -- ADDR 1696
			"00000000000000000000000000000000" , -- ADDR 1697
			"00000000000000000000000000000000" , -- ADDR 1698
			"00000000000000000000000000000000" , -- ADDR 1699
			"00000000000000000000000000000000" , -- ADDR 1700
			"00000000000000000000000000000000" , -- ADDR 1701
			"00000000000000000000000000000000" , -- ADDR 1702
			"00000000000000000000000000000000" , -- ADDR 1703
			"00000000000000000000000000000000" , -- ADDR 1704
			"00000000000000000000000000000000" , -- ADDR 1705
			"00000000000000000000000000000000" , -- ADDR 1706
			"00000000000000000000000000000000" , -- ADDR 1707
			"00000000000000000000000000000000" , -- ADDR 1708
			"00000000000000000000000000000000" , -- ADDR 1709
			"00000000000000000000000000000000" , -- ADDR 1710
			"00000000000000000000000000000000" , -- ADDR 1711
			"00000000000000000000000000000000" , -- ADDR 1712
			"00000000000000000000000000000000" , -- ADDR 1713
			"00000000000000000000000000000000" , -- ADDR 1714
			"00000000000000000000000000000000" , -- ADDR 1715
			"00000000000000000000000000000000" , -- ADDR 1716
			"00000000000000000000000000000000" , -- ADDR 1717
			"00000000000000000000000000000000" , -- ADDR 1718
			"00000000000000000000000000000000" , -- ADDR 1719
			"00000000000000000000000000000000" , -- ADDR 1720
			"00000000000000000000000000000000" , -- ADDR 1721
			"00000000000000000000000000000000" , -- ADDR 1722
			"00000000000000000000000000000000" , -- ADDR 1723
			"00000000000000000000000000000000" , -- ADDR 1724
			"00000000000000000000000000000000" , -- ADDR 1725
			"00000000000000000000000000000000" , -- ADDR 1726
			"00000000000000000000000000000000" , -- ADDR 1727
			"00000000000000000000000000000000" , -- ADDR 1728
			"00000000000000000000000000000000" , -- ADDR 1729
			"00000000000000000000000000000000" , -- ADDR 1730
			"00000000000000000000000000000000" , -- ADDR 1731
			"00000000000000000000000000000000" , -- ADDR 1732
			"00000000000000000000000000000000" , -- ADDR 1733
			"00000000000000000000000000000000" , -- ADDR 1734
			"00000000000000000000000000000000" , -- ADDR 1735
			"00000000000000000000000000000000" , -- ADDR 1736
			"00000000000000000000000000000000" , -- ADDR 1737
			"00000000000000000000000000000000" , -- ADDR 1738
			"00000000000000000000000000000000" , -- ADDR 1739
			"00000000000000000000000000000000" , -- ADDR 1740
			"00000000000000000000000000000000" , -- ADDR 1741
			"00000000000000000000000000000000" , -- ADDR 1742
			"00000000000000000000000000000000" , -- ADDR 1743
			"00000000000000000000000000000000" , -- ADDR 1744
			"00000000000000000000000000000000" , -- ADDR 1745
			"00000000000000000000000000000000" , -- ADDR 1746
			"00000000000000000000000000000000" , -- ADDR 1747
			"00000000000000000000000000000000" , -- ADDR 1748
			"00000000000000000000000000000000" , -- ADDR 1749
			"00000000000000000000000000000000" , -- ADDR 1750
			"00000000000000000000000000000000" , -- ADDR 1751
			"00000000000000000000000000000000" , -- ADDR 1752
			"00000000000000000000000000000000" , -- ADDR 1753
			"00000000000000000000000000000000" , -- ADDR 1754
			"00000000000000000000000000000000" , -- ADDR 1755
			"00000000000000000000000000000000" , -- ADDR 1756
			"00000000000000000000000000000000" , -- ADDR 1757
			"00000000000000000000000000000000" , -- ADDR 1758
			"00000000000000000000000000000000" , -- ADDR 1759
			"00000000000000000000000000000000" , -- ADDR 1760
			"00000000000000000000000000000000" , -- ADDR 1761
			"00000000000000000000000000000000" , -- ADDR 1762
			"00000000000000000000000000000000" , -- ADDR 1763
			"00000000000000000000000000000000" , -- ADDR 1764
			"00000000000000000000000000000000" , -- ADDR 1765
			"00000000000000000000000000000000" , -- ADDR 1766
			"00000000000000000000000000000000" , -- ADDR 1767
			"00000000000000000000000000000000" , -- ADDR 1768
			"00000000000000000000000000000000" , -- ADDR 1769
			"00000000000000000000000000000000" , -- ADDR 1770
			"00000000000000000000000000000000" , -- ADDR 1771
			"00000000000000000000000000000000" , -- ADDR 1772
			"00000000000000000000000000000000" , -- ADDR 1773
			"00000000000000000000000000000000" , -- ADDR 1774
			"00000000000000000000000000000000" , -- ADDR 1775
			"00000000000000000000000000000000" , -- ADDR 1776
			"00000000000000000000000000000000" , -- ADDR 1777
			"00000000000000000000000000000000" , -- ADDR 1778
			"00000000000000000000000000000000" , -- ADDR 1779
			"00000000000000000000000000000000" , -- ADDR 1780
			"00000000000000000000000000000000" , -- ADDR 1781
			"00000000000000000000000000000000" , -- ADDR 1782
			"00000000000000000000000000000000" , -- ADDR 1783
			"00000000000000000000000000000000" , -- ADDR 1784
			"00000000000000000000000000000000" , -- ADDR 1785
			"00000000000000000000000000000000" , -- ADDR 1786
			"00000000000000000000000000000000" , -- ADDR 1787
			"00000000000000000000000000000000" , -- ADDR 1788
			"00000000000000000000000000000000" , -- ADDR 1789
			"00000000000000000000000000000000" , -- ADDR 1790
			"00000000000000000000000000000000" , -- ADDR 1791
			"00000000000000000000000000000000" , -- ADDR 1792
			"00000000000000000000000000000000" , -- ADDR 1793
			"00000000000000000000000000000000" , -- ADDR 1794
			"00000000000000000000000000000000" , -- ADDR 1795
			"00000000000000000000000000000000" , -- ADDR 1796
			"00000000000000000000000000000000" , -- ADDR 1797
			"00000000000000000000000000000000" , -- ADDR 1798
			"00000000000000000000000000000000" , -- ADDR 1799
			"00000000000000000000000000000000" , -- ADDR 1800
			"00000000000000000000000000000000" , -- ADDR 1801
			"00000000000000000000000000000000" , -- ADDR 1802
			"00000000000000000000000000000000" , -- ADDR 1803
			"00000000000000000000000000000000" , -- ADDR 1804
			"00000000000000000000000000000000" , -- ADDR 1805
			"00000000000000000000000000000000" , -- ADDR 1806
			"00000000000000000000000000000000" , -- ADDR 1807
			"00000000000000000000000000000000" , -- ADDR 1808
			"00000000000000000000000000000000" , -- ADDR 1809
			"00000000000000000000000000000000" , -- ADDR 1810
			"00000000000000000000000000000000" , -- ADDR 1811
			"00000000000000000000000000000000" , -- ADDR 1812
			"00000000000000000000000000000000" , -- ADDR 1813
			"00000000000000000000000000000000" , -- ADDR 1814
			"00000000000000000000000000000000" , -- ADDR 1815
			"00000000000000000000000000000000" , -- ADDR 1816
			"00000000000000000000000000000000" , -- ADDR 1817
			"00000000000000000000000000000000" , -- ADDR 1818
			"00000000000000000000000000000000" , -- ADDR 1819
			"00000000000000000000000000000000" , -- ADDR 1820
			"00000000000000000000000000000000" , -- ADDR 1821
			"00000000000000000000000000000000" , -- ADDR 1822
			"00000000000000000000000000000000" , -- ADDR 1823
			"00000000000000000000000000000000" , -- ADDR 1824
			"00000000000000000000000000000000" , -- ADDR 1825
			"00000000000000000000000000000000" , -- ADDR 1826
			"00000000000000000000000000000000" , -- ADDR 1827
			"00000000000000000000000000000000" , -- ADDR 1828
			"00000000000000000000000000000000" , -- ADDR 1829
			"00000000000000000000000000000000" , -- ADDR 1830
			"00000000000000000000000000000000" , -- ADDR 1831
			"00000000000000000000000000000000" , -- ADDR 1832
			"00000000000000000000000000000000" , -- ADDR 1833
			"00000000000000000000000000000000" , -- ADDR 1834
			"00000000000000000000000000000000" , -- ADDR 1835
			"00000000000000000000000000000000" , -- ADDR 1836
			"00000000000000000000000000000000" , -- ADDR 1837
			"00000000000000000000000000000000" , -- ADDR 1838
			"00000000000000000000000000000000" , -- ADDR 1839
			"00000000000000000000000000000000" , -- ADDR 1840
			"00000000000000000000000000000000" , -- ADDR 1841
			"00000000000000000000000000000000" , -- ADDR 1842
			"00000000000000000000000000000000" , -- ADDR 1843
			"00000000000000000000000000000000" , -- ADDR 1844
			"00000000000000000000000000000000" , -- ADDR 1845
			"00000000000000000000000000000000" , -- ADDR 1846
			"00000000000000000000000000000000" , -- ADDR 1847
			"00000000000000000000000000000000" , -- ADDR 1848
			"00000000000000000000000000000000" , -- ADDR 1849
			"00000000000000000000000000000000" , -- ADDR 1850
			"00000000000000000000000000000000" , -- ADDR 1851
			"00000000000000000000000000000000" , -- ADDR 1852
			"00000000000000000000000000000000" , -- ADDR 1853
			"00000000000000000000000000000000" , -- ADDR 1854
			"00000000000000000000000000000000" , -- ADDR 1855
			"00000000000000000000000000000000" , -- ADDR 1856
			"00000000000000000000000000000000" , -- ADDR 1857
			"00000000000000000000000000000000" , -- ADDR 1858
			"00000000000000000000000000000000" , -- ADDR 1859
			"00000000000000000000000000000000" , -- ADDR 1860
			"00000000000000000000000000000000" , -- ADDR 1861
			"00000000000000000000000000000000" , -- ADDR 1862
			"00000000000000000000000000000000" , -- ADDR 1863
			"00000000000000000000000000000000" , -- ADDR 1864
			"00000000000000000000000000000000" , -- ADDR 1865
			"00000000000000000000000000000000" , -- ADDR 1866
			"00000000000000000000000000000000" , -- ADDR 1867
			"00000000000000000000000000000000" , -- ADDR 1868
			"00000000000000000000000000000000" , -- ADDR 1869
			"00000000000000000000000000000000" , -- ADDR 1870
			"00000000000000000000000000000000" , -- ADDR 1871
			"00000000000000000000000000000000" , -- ADDR 1872
			"00000000000000000000000000000000" , -- ADDR 1873
			"00000000000000000000000000000000" , -- ADDR 1874
			"00000000000000000000000000000000" , -- ADDR 1875
			"00000000000000000000000000000000" , -- ADDR 1876
			"00000000000000000000000000000000" , -- ADDR 1877
			"00000000000000000000000000000000" , -- ADDR 1878
			"00000000000000000000000000000000" , -- ADDR 1879
			"00000000000000000000000000000000" , -- ADDR 1880
			"00000000000000000000000000000000" , -- ADDR 1881
			"00000000000000000000000000000000" , -- ADDR 1882
			"00000000000000000000000000000000" , -- ADDR 1883
			"00000000000000000000000000000000" , -- ADDR 1884
			"00000000000000000000000000000000" , -- ADDR 1885
			"00000000000000000000000000000000" , -- ADDR 1886
			"00000000000000000000000000000000" , -- ADDR 1887
			"00000000000000000000000000000000" , -- ADDR 1888
			"00000000000000000000000000000000" , -- ADDR 1889
			"00000000000000000000000000000000" , -- ADDR 1890
			"00000000000000000000000000000000" , -- ADDR 1891
			"00000000000000000000000000000000" , -- ADDR 1892
			"00000000000000000000000000000000" , -- ADDR 1893
			"00000000000000000000000000000000" , -- ADDR 1894
			"00000000000000000000000000000000" , -- ADDR 1895
			"00000000000000000000000000000000" , -- ADDR 1896
			"00000000000000000000000000000000" , -- ADDR 1897
			"00000000000000000000000000000000" , -- ADDR 1898
			"00000000000000000000000000000000" , -- ADDR 1899
			"00000000000000000000000000000000" , -- ADDR 1900
			"00000000000000000000000000000000" , -- ADDR 1901
			"00000000000000000000000000000000" , -- ADDR 1902
			"00000000000000000000000000000000" , -- ADDR 1903
			"00000000000000000000000000000000" , -- ADDR 1904
			"00000000000000000000000000000000" , -- ADDR 1905
			"00000000000000000000000000000000" , -- ADDR 1906
			"00000000000000000000000000000000" , -- ADDR 1907
			"00000000000000000000000000000000" , -- ADDR 1908
			"00000000000000000000000000000000" , -- ADDR 1909
			"00000000000000000000000000000000" , -- ADDR 1910
			"00000000000000000000000000000000" , -- ADDR 1911
			"00000000000000000000000000000000" , -- ADDR 1912
			"00000000000000000000000000000000" , -- ADDR 1913
			"00000000000000000000000000000000" , -- ADDR 1914
			"00000000000000000000000000000000" , -- ADDR 1915
			"00000000000000000000000000000000" , -- ADDR 1916
			"00000000000000000000000000000000" , -- ADDR 1917
			"00000000000000000000000000000000" , -- ADDR 1918
			"00000000000000000000000000000000" , -- ADDR 1919
			"00000000000000000000000000000000" , -- ADDR 1920
			"00000000000000000000000000000000" , -- ADDR 1921
			"00000000000000000000000000000000" , -- ADDR 1922
			"00000000000000000000000000000000" , -- ADDR 1923
			"00000000000000000000000000000000" , -- ADDR 1924
			"00000000000000000000000000000000" , -- ADDR 1925
			"00000000000000000000000000000000" , -- ADDR 1926
			"00000000000000000000000000000000" , -- ADDR 1927
			"00000000000000000000000000000000" , -- ADDR 1928
			"00000000000000000000000000000000" , -- ADDR 1929
			"00000000000000000000000000000000" , -- ADDR 1930
			"00000000000000000000000000000000" , -- ADDR 1931
			"00000000000000000000000000000000" , -- ADDR 1932
			"00000000000000000000000000000000" , -- ADDR 1933
			"00000000000000000000000000000000" , -- ADDR 1934
			"00000000000000000000000000000000" , -- ADDR 1935
			"00000000000000000000000000000000" , -- ADDR 1936
			"00000000000000000000000000000000" , -- ADDR 1937
			"00000000000000000000000000000000" , -- ADDR 1938
			"00000000000000000000000000000000" , -- ADDR 1939
			"00000000000000000000000000000000" , -- ADDR 1940
			"00000000000000000000000000000000" , -- ADDR 1941
			"00000000000000000000000000000000" , -- ADDR 1942
			"00000000000000000000000000000000" , -- ADDR 1943
			"00000000000000000000000000000000" , -- ADDR 1944
			"00000000000000000000000000000000" , -- ADDR 1945
			"00000000000000000000000000000000" , -- ADDR 1946
			"00000000000000000000000000000000" , -- ADDR 1947
			"00000000000000000000000000000000" , -- ADDR 1948
			"00000000000000000000000000000000" , -- ADDR 1949
			"00000000000000000000000000000000" , -- ADDR 1950
			"00000000000000000000000000000000" , -- ADDR 1951
			"00000000000000000000000000000000" , -- ADDR 1952
			"00000000000000000000000000000000" , -- ADDR 1953
			"00000000000000000000000000000000" , -- ADDR 1954
			"00000000000000000000000000000000" , -- ADDR 1955
			"00000000000000000000000000000000" , -- ADDR 1956
			"00000000000000000000000000000000" , -- ADDR 1957
			"00000000000000000000000000000000" , -- ADDR 1958
			"00000000000000000000000000000000" , -- ADDR 1959
			"00000000000000000000000000000000" , -- ADDR 1960
			"00000000000000000000000000000000" , -- ADDR 1961
			"00000000000000000000000000000000" , -- ADDR 1962
			"00000000000000000000000000000000" , -- ADDR 1963
			"00000000000000000000000000000000" , -- ADDR 1964
			"00000000000000000000000000000000" , -- ADDR 1965
			"00000000000000000000000000000000" , -- ADDR 1966
			"00000000000000000000000000000000" , -- ADDR 1967
			"00000000000000000000000000000000" , -- ADDR 1968
			"00000000000000000000000000000000" , -- ADDR 1969
			"00000000000000000000000000000000" , -- ADDR 1970
			"00000000000000000000000000000000" , -- ADDR 1971
			"00000000000000000000000000000000" , -- ADDR 1972
			"00000000000000000000000000000000" , -- ADDR 1973
			"00000000000000000000000000000000" , -- ADDR 1974
			"00000000000000000000000000000000" , -- ADDR 1975
			"00000000000000000000000000000000" , -- ADDR 1976
			"00000000000000000000000000000000" , -- ADDR 1977
			"00000000000000000000000000000000" , -- ADDR 1978
			"00000000000000000000000000000000" , -- ADDR 1979
			"00000000000000000000000000000000" , -- ADDR 1980
			"00000000000000000000000000000000" , -- ADDR 1981
			"00000000000000000000000000000000" , -- ADDR 1982
			"00000000000000000000000000000000" , -- ADDR 1983
			"00000000000000000000000000000000" , -- ADDR 1984
			"00000000000000000000000000000000" , -- ADDR 1985
			"00000000000000000000000000000000" , -- ADDR 1986
			"00000000000000000000000000000000" , -- ADDR 1987
			"00000000000000000000000000000000" , -- ADDR 1988
			"00000000000000000000000000000000" , -- ADDR 1989
			"00000000000000000000000000000000" , -- ADDR 1990
			"00000000000000000000000000000000" , -- ADDR 1991
			"00000000000000000000000000000000" , -- ADDR 1992
			"00000000000000000000000000000000" , -- ADDR 1993
			"00000000000000000000000000000000" , -- ADDR 1994
			"00000000000000000000000000000000" , -- ADDR 1995
			"00000000000000000000000000000000" , -- ADDR 1996
			"00000000000000000000000000000000" , -- ADDR 1997
			"00000000000000000000000000000000" , -- ADDR 1998
			"00000000000000000000000000000000" , -- ADDR 1999
			"00000000000000000000000000000000" , -- ADDR 2000
			"00000000000000000000000000000000" , -- ADDR 2001
			"00000000000000000000000000000000" , -- ADDR 2002
			"00000000000000000000000000000000" , -- ADDR 2003
			"00000000000000000000000000000000" , -- ADDR 2004
			"00000000000000000000000000000000" , -- ADDR 2005
			"00000000000000000000000000000000" , -- ADDR 2006
			"00000000000000000000000000000000" , -- ADDR 2007
			"00000000000000000000000000000000" , -- ADDR 2008
			"00000000000000000000000000000000" , -- ADDR 2009
			"00000000000000000000000000000000" , -- ADDR 2010
			"00000000000000000000000000000000" , -- ADDR 2011
			"00000000000000000000000000000000" , -- ADDR 2012
			"00000000000000000000000000000000" , -- ADDR 2013
			"00000000000000000000000000000000" , -- ADDR 2014
			"00000000000000000000000000000000" , -- ADDR 2015
			"00000000000000000000000000000000" , -- ADDR 2016
			"00000000000000000000000000000000" , -- ADDR 2017
			"00000000000000000000000000000000" , -- ADDR 2018
			"00000000000000000000000000000000" , -- ADDR 2019
			"00000000000000000000000000000000" , -- ADDR 2020
			"00000000000000000000000000000000" , -- ADDR 2021
			"00000000000000000000000000000000" , -- ADDR 2022
			"00000000000000000000000000000000" , -- ADDR 2023
			"00000000000000000000000000000000" , -- ADDR 2024
			"00000000000000000000000000000000" , -- ADDR 2025
			"00000000000000000000000000000000" , -- ADDR 2026
			"00000000000000000000000000000000" , -- ADDR 2027
			"00000000000000000000000000000000" , -- ADDR 2028
			"00000000000000000000000000000000" , -- ADDR 2029
			"00000000000000000000000000000000" , -- ADDR 2030
			"00000000000000000000000000000000" , -- ADDR 2031
			"00000000000000000000000000000000" , -- ADDR 2032
			"00000000000000000000000000000000" , -- ADDR 2033
			"00000000000000000000000000000000" , -- ADDR 2034
			"00000000000000000000000000000000" , -- ADDR 2035
			"00000000000000000000000000000000" , -- ADDR 2036
			"00000000000000000000000000000000" , -- ADDR 2037
			"00000000000000000000000000000000" , -- ADDR 2038
			"00000000000000000000000000000000" , -- ADDR 2039
			"00000000000000000000000000000000" , -- ADDR 2040
			"00000000000000000000000000000000" , -- ADDR 2041
			"00000000000000000000000000000000" , -- ADDR 2042
			"00000000000000000000000000000000" , -- ADDR 2043
			"00000000000000000000000000000000" , -- ADDR 2044
			"00000000000000000000000000000000" , -- ADDR 2045
			"00000000000000000000000000000000" , -- ADDR 2046
			"00000000000000000000000000000000"   -- ADDR 2047
			);
			
begin
	
	process (CLK)
	begin
		if (rising_edge(CLK)) then
			-- In the case of Altera Quartus, it is extremely essential that the output assignment stays in the process.
			-- Otherwise, Altera Quartus will not infer the VHDL code as ROM.
			-- However, in the case of Xilinx ISE, it does not matter whether the output assignment stays in the process
			-- or outside of it with synchronization to the clock pulse by another signal. The VHDL code will infer as ROM anyway.
			DATA <= ROM (to_integer(unsigned(ADDR)));
		end if;
	end process;
	
end Behavioral;

-- Extremely important: In order for Altera Quartus to infer the VHDL code as ROM, the setting in the path
-- "Assignments/Device…/Device and Pin Options…/Configuration/Configuration mode" must be changed to
-- "Single Uncompressed Image with memory initialization (512 Kbits UFM)".

