----------------------------------------------------------------------------------------------------
-- Author           : Pourya Khodagholipour (P.KH)
-- Project Name     : HBA (Hardware Bee Algorithm)
-- File Name        : TSP_Y_One_Port_ROM_Sync
-- Module Name      : TSP_Y_One_Port_ROM_Sync
-- HDL Standard     : VHDL
-- Approach         : Behavioral
-- Description      : Single-port ROM with synchronous read (Block RAM)
-- Comments         : eil51 Database Y Coordinates
-- Dependencies     : ---
-- Target Devices   : Virtex 5 - XC5VLX330
-- Speed Estimation : ---
-- Area  Estimation : 1 RAM/FIFO
-- Tools            : ISE Design Suite v14.7 - Altera Quartus 16.1 Lite
-- Module Version   : 
-- Creation Date    : 2016/08
-- Revision Date    : 2024/07/10
----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity TSP_Y_One_Port_ROM_Sync is
	generic (
				ADDR_WIDTH : natural := 8;
				DATA_WIDTH : natural := 24);
	port    (
				CLK        : in  std_logic;
				ADDR       : in  std_logic_vector (ADDR_WIDTH-1 downto 0);
				DATA       : out std_logic_vector (DATA_WIDTH-1 downto 0));
end TSP_Y_One_Port_ROM_Sync;

architecture Behavioral of TSP_Y_One_Port_ROM_Sync is
	
	type ROM_Type is array (0 to 2**ADDR_WIDTH-1) of STD_LOGIC_VECTOR (DATA_WIDTH-1 downto 0);
	constant ROM : ROM_Type := (
		"000000001100101100100000" , -- ADDR 0
		"000000001011111101101000" , -- ADDR 1
		"000000001111101000000000" , -- ADDR 2
		"000000000110010110010000" , -- ADDR 3
		"000000000111010100110000" , -- ADDR 4
		"000000001011011110011000" , -- ADDR 5
		"000000001111011000011000" , -- ADDR 6
		"000000001111001000110000" , -- ADDR 7
		"000000001000000011101000" , -- ADDR 8
		"000000000101001000001000" , -- ADDR 9
		"000000001010000000101000" , -- ADDR 10
		"000000000111110100000000" , -- ADDR 11
		"000000000110000110101000" , -- ADDR 12
		"000000001010010000010000" , -- ADDR 13
		"000000000011111010000000" , -- ADDR 14
		"000000001010000000101000" , -- ADDR 15
		"000000000101100111011000" , -- ADDR 16
		"000000001000000011101000" , -- ADDR 17
		"000000000011001011001000" , -- ADDR 18
		"000000001110001010010000" , -- ADDR 19
		"000000001010010000010000" , -- ADDR 20
		"000000001101111010101000" , -- ADDR 21
		"000000001101111010101000" , -- ADDR 22
		"000000001100101100100000" , -- ADDR 23
		"000000001001010001110000" , -- ADDR 24
		"000000010000100110100000" , -- ADDR 25
		"000000001011101110000000" , -- ADDR 26
		"000000010000010110111000" , -- ADDR 27
		"000000001011101110000000" , -- ADDR 28
		"000000000110100101111000" , -- ADDR 29
		"000000010000110110001000" , -- ADDR 30
		"000000001011001110110000" , -- ADDR 31
		"000000000010011100010000" , -- ADDR 32
		"000000001000000011101000" , -- ADDR 33
		"000000001111011000011000" , -- ADDR 34
		"000000010000110110001000" , -- ADDR 35
		"000000000101010111110000" , -- ADDR 36
		"000000001000100010111000" , -- ADDR 37
		"000000000011101010011000" , -- ADDR 38
		"000000000001011101110000" , -- ADDR 39
		"000000000100001001101000" , -- ADDR 40
		"000000000010011100010000" , -- ADDR 41
		"000000001111101000000000" , -- ADDR 42
		"000000000011101010011000" , -- ADDR 43
		"000000000010011100010000" , -- ADDR 44
		"000000001001100001011000" , -- ADDR 45
		"000000000111110100000000" , -- ADDR 46
		"000000001101011011011000" , -- ADDR 47
		"000000000110110101100000" , -- ADDR 48
		"000000001001000010001000" , -- ADDR 49
		"000000001001110001000000" , -- ADDR 50
		"000000000000000000000000" , -- ADDR 51
		"000000000000000000000000" , -- ADDR 52
		"000000000000000000000000" , -- ADDR 53
		"000000000000000000000000" , -- ADDR 54
		"000000000000000000000000" , -- ADDR 55
		"000000000000000000000000" , -- ADDR 56
		"000000000000000000000000" , -- ADDR 57
		"000000000000000000000000" , -- ADDR 58
		"000000000000000000000000" , -- ADDR 59
		"000000000000000000000000" , -- ADDR 60
		"000000000000000000000000" , -- ADDR 61
		"000000000000000000000000" , -- ADDR 62
		"000000000000000000000000" , -- ADDR 63
		"000000000000000000000000" , -- ADDR 64
		"000000000000000000000000" , -- ADDR 65
		"000000000000000000000000" , -- ADDR 66
		"000000000000000000000000" , -- ADDR 67
		"000000000000000000000000" , -- ADDR 68
		"000000000000000000000000" , -- ADDR 69
		"000000000000000000000000" , -- ADDR 70
		"000000000000000000000000" , -- ADDR 71
		"000000000000000000000000" , -- ADDR 72
		"000000000000000000000000" , -- ADDR 73
		"000000000000000000000000" , -- ADDR 74
		"000000000000000000000000" , -- ADDR 75
		"000000000000000000000000" , -- ADDR 76
		"000000000000000000000000" , -- ADDR 77
		"000000000000000000000000" , -- ADDR 78
		"000000000000000000000000" , -- ADDR 79
		"000000000000000000000000" , -- ADDR 80
		"000000000000000000000000" , -- ADDR 81
		"000000000000000000000000" , -- ADDR 82
		"000000000000000000000000" , -- ADDR 83
		"000000000000000000000000" , -- ADDR 84
		"000000000000000000000000" , -- ADDR 85
		"000000000000000000000000" , -- ADDR 86
		"000000000000000000000000" , -- ADDR 87
		"000000000000000000000000" , -- ADDR 88
		"000000000000000000000000" , -- ADDR 89
		"000000000000000000000000" , -- ADDR 90
		"000000000000000000000000" , -- ADDR 91
		"000000000000000000000000" , -- ADDR 92
		"000000000000000000000000" , -- ADDR 93
		"000000000000000000000000" , -- ADDR 94
		"000000000000000000000000" , -- ADDR 95
		"000000000000000000000000" , -- ADDR 96
		"000000000000000000000000" , -- ADDR 97
		"000000000000000000000000" , -- ADDR 98
		"000000000000000000000000" , -- ADDR 99
		"000000000000000000000000" , -- ADDR 100
		"000000000000000000000000" , -- ADDR 101
		"000000000000000000000000" , -- ADDR 102
		"000000000000000000000000" , -- ADDR 103
		"000000000000000000000000" , -- ADDR 104
		"000000000000000000000000" , -- ADDR 105
		"000000000000000000000000" , -- ADDR 106
		"000000000000000000000000" , -- ADDR 107
		"000000000000000000000000" , -- ADDR 108
		"000000000000000000000000" , -- ADDR 109
		"000000000000000000000000" , -- ADDR 110
		"000000000000000000000000" , -- ADDR 111
		"000000000000000000000000" , -- ADDR 112
		"000000000000000000000000" , -- ADDR 113
		"000000000000000000000000" , -- ADDR 114
		"000000000000000000000000" , -- ADDR 115
		"000000000000000000000000" , -- ADDR 116
		"000000000000000000000000" , -- ADDR 117
		"000000000000000000000000" , -- ADDR 118
		"000000000000000000000000" , -- ADDR 119
		"000000000000000000000000" , -- ADDR 120
		"000000000000000000000000" , -- ADDR 121
		"000000000000000000000000" , -- ADDR 122
		"000000000000000000000000" , -- ADDR 123
		"000000000000000000000000" , -- ADDR 124
		"000000000000000000000000" , -- ADDR 125
		"000000000000000000000000" , -- ADDR 126
		"000000000000000000000000" , -- ADDR 127
		"000000000000000000000000" , -- ADDR 128
		"000000000000000000000000" , -- ADDR 129
		"000000000000000000000000" , -- ADDR 130
		"000000000000000000000000" , -- ADDR 131
		"000000000000000000000000" , -- ADDR 132
		"000000000000000000000000" , -- ADDR 133
		"000000000000000000000000" , -- ADDR 134
		"000000000000000000000000" , -- ADDR 135
		"000000000000000000000000" , -- ADDR 136
		"000000000000000000000000" , -- ADDR 137
		"000000000000000000000000" , -- ADDR 138
		"000000000000000000000000" , -- ADDR 139
		"000000000000000000000000" , -- ADDR 140
		"000000000000000000000000" , -- ADDR 141
		"000000000000000000000000" , -- ADDR 142
		"000000000000000000000000" , -- ADDR 143
		"000000000000000000000000" , -- ADDR 144
		"000000000000000000000000" , -- ADDR 145
		"000000000000000000000000" , -- ADDR 146
		"000000000000000000000000" , -- ADDR 147
		"000000000000000000000000" , -- ADDR 148
		"000000000000000000000000" , -- ADDR 149
		"000000000000000000000000" , -- ADDR 150
		"000000000000000000000000" , -- ADDR 151
		"000000000000000000000000" , -- ADDR 152
		"000000000000000000000000" , -- ADDR 153
		"000000000000000000000000" , -- ADDR 154
		"000000000000000000000000" , -- ADDR 155
		"000000000000000000000000" , -- ADDR 156
		"000000000000000000000000" , -- ADDR 157
		"000000000000000000000000" , -- ADDR 158
		"000000000000000000000000" , -- ADDR 159
		"000000000000000000000000" , -- ADDR 160
		"000000000000000000000000" , -- ADDR 161
		"000000000000000000000000" , -- ADDR 162
		"000000000000000000000000" , -- ADDR 163
		"000000000000000000000000" , -- ADDR 164
		"000000000000000000000000" , -- ADDR 165
		"000000000000000000000000" , -- ADDR 166
		"000000000000000000000000" , -- ADDR 167
		"000000000000000000000000" , -- ADDR 168
		"000000000000000000000000" , -- ADDR 169
		"000000000000000000000000" , -- ADDR 170
		"000000000000000000000000" , -- ADDR 171
		"000000000000000000000000" , -- ADDR 172
		"000000000000000000000000" , -- ADDR 173
		"000000000000000000000000" , -- ADDR 174
		"000000000000000000000000" , -- ADDR 175
		"000000000000000000000000" , -- ADDR 176
		"000000000000000000000000" , -- ADDR 177
		"000000000000000000000000" , -- ADDR 178
		"000000000000000000000000" , -- ADDR 179
		"000000000000000000000000" , -- ADDR 180
		"000000000000000000000000" , -- ADDR 181
		"000000000000000000000000" , -- ADDR 182
		"000000000000000000000000" , -- ADDR 183
		"000000000000000000000000" , -- ADDR 184
		"000000000000000000000000" , -- ADDR 185
		"000000000000000000000000" , -- ADDR 186
		"000000000000000000000000" , -- ADDR 187
		"000000000000000000000000" , -- ADDR 188
		"000000000000000000000000" , -- ADDR 189
		"000000000000000000000000" , -- ADDR 190
		"000000000000000000000000" , -- ADDR 191
		"000000000000000000000000" , -- ADDR 192
		"000000000000000000000000" , -- ADDR 193
		"000000000000000000000000" , -- ADDR 194
		"000000000000000000000000" , -- ADDR 195
		"000000000000000000000000" , -- ADDR 196
		"000000000000000000000000" , -- ADDR 197
		"000000000000000000000000" , -- ADDR 198
		"000000000000000000000000" , -- ADDR 199
		"000000000000000000000000" , -- ADDR 200
		"000000000000000000000000" , -- ADDR 201
		"000000000000000000000000" , -- ADDR 202
		"000000000000000000000000" , -- ADDR 203
		"000000000000000000000000" , -- ADDR 204
		"000000000000000000000000" , -- ADDR 205
		"000000000000000000000000" , -- ADDR 206
		"000000000000000000000000" , -- ADDR 207
		"000000000000000000000000" , -- ADDR 208
		"000000000000000000000000" , -- ADDR 209
		"000000000000000000000000" , -- ADDR 210
		"000000000000000000000000" , -- ADDR 211
		"000000000000000000000000" , -- ADDR 212
		"000000000000000000000000" , -- ADDR 213
		"000000000000000000000000" , -- ADDR 214
		"000000000000000000000000" , -- ADDR 215
		"000000000000000000000000" , -- ADDR 216
		"000000000000000000000000" , -- ADDR 217
		"000000000000000000000000" , -- ADDR 218
		"000000000000000000000000" , -- ADDR 219
		"000000000000000000000000" , -- ADDR 220
		"000000000000000000000000" , -- ADDR 221
		"000000000000000000000000" , -- ADDR 222
		"000000000000000000000000" , -- ADDR 223
		"000000000000000000000000" , -- ADDR 224
		"000000000000000000000000" , -- ADDR 225
		"000000000000000000000000" , -- ADDR 226
		"000000000000000000000000" , -- ADDR 227
		"000000000000000000000000" , -- ADDR 228
		"000000000000000000000000" , -- ADDR 229
		"000000000000000000000000" , -- ADDR 230
		"000000000000000000000000" , -- ADDR 231
		"000000000000000000000000" , -- ADDR 232
		"000000000000000000000000" , -- ADDR 233
		"000000000000000000000000" , -- ADDR 234
		"000000000000000000000000" , -- ADDR 235
		"000000000000000000000000" , -- ADDR 236
		"000000000000000000000000" , -- ADDR 237
		"000000000000000000000000" , -- ADDR 238
		"000000000000000000000000" , -- ADDR 239
		"000000000000000000000000" , -- ADDR 240
		"000000000000000000000000" , -- ADDR 241
		"000000000000000000000000" , -- ADDR 242
		"000000000000000000000000" , -- ADDR 243
		"000000000000000000000000" , -- ADDR 244
		"000000000000000000000000" , -- ADDR 245
		"000000000000000000000000" , -- ADDR 246
		"000000000000000000000000" , -- ADDR 247
		"000000000000000000000000" , -- ADDR 248
		"000000000000000000000000" , -- ADDR 249
		"000000000000000000000000" , -- ADDR 250
		"000000000000000000000000" , -- ADDR 251
		"000000000000000000000000" , -- ADDR 252
		"000000000000000000000000" , -- ADDR 253
		"000000000000000000000000" , -- ADDR 254
		"000000000000000000000000"   -- ADDR 255
	);
			
begin
	
	process (CLK)
	begin
		if (rising_edge(CLK)) then
			-- In the case of Altera Quartus, it is extremely essential that the output assignment stays in the process.
			-- Otherwise, Altera Quartus will not infer the VHDL code as ROM.
			-- However, in the case of Xilinx ISE, it does not matter whether the output assignment stays in the process
			-- or outside of it with synchronization to the clock pulse by another signal. The VHDL code will infer as ROM anyway.
			DATA <= ROM (to_integer(unsigned(ADDR)));
		end if;
	end process;
	
end Behavioral;

-- Extremely important: In order for Altera Quartus to infer the VHDL code as ROM, the setting in the path
-- "Assignments/Device…/Device and Pin Options…/Configuration/Configuration mode" must be changed to
-- "Single Uncompressed Image with memory initialization (512 Kbits UFM)".