----------------------------------------------------------------------------------------------------
-- Author           : Pourya Khodagholipour (P.KH)
-- Project Name     : HBA (Hardware Bee Algorithm)
-- File Name        : TSP_Dist_One_Port_ROM_Sync
-- Module Name      : TSP_Dist_One_Port_ROM_Sync
-- HDL Standard     : VHDL
-- Approach         : Behavioral
-- Description      : Single-port ROM with synchronous read (Block RAM)
-- Comments         : eil51 Database Distance matrix
-- Dependencies     : ---
-- Target Devices   : Virtex 5 - XC5VLX330
-- Speed Estimation : ---
-- Area  Estimation : 2 RAM/FIFO
-- Tools            : ISE Design Suite v14.7 - Altera Quartus 16.1 Lite
-- Module Version   : 
-- Creation Date    : 2016/08
-- Revision Date    : 2024/07/08
----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity TSP_Dist_One_Port_ROM_Sync is
	generic (
				ADDR_WIDTH : natural := 11;
				DATA_WIDTH : natural := 32);
	port    (
				CLK        : in  std_logic;
				ADDR       : in  std_logic_vector (ADDR_WIDTH-1 downto 0);
				DATA       : out std_logic_vector (DATA_WIDTH-1 downto 0));
end TSP_Dist_One_Port_ROM_Sync;

architecture Behavioral of TSP_Dist_One_Port_ROM_Sync is

	type ROM_Type is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector (DATA_WIDTH-1 downto 0);
	constant ROM : ROM_Type := (
			"11111111111111111111111111111111" , -- ADDR 0
			"00000000000000000011000001010001" , -- ADDR 1
			"00000000000000000100101100001001" , -- ADDR 2
			"00000000000000000111100101011000" , -- ADDR 3
			"00000000000000000101011010111100" , -- ADDR 4
			"00000000000000000100000101111011" , -- ADDR 5
			"00000000000000000101100100101001" , -- ADDR 6
			"00000000000000000010110110001110" , -- ADDR 7
			"00000000000000000101111010001111" , -- ADDR 8
			"00000000000000001000010011011111" , -- ADDR 9
			"00000000000000000010111100110011" , -- ADDR 10
			"00000000000000000101000110010001" , -- ADDR 11
			"00000000000000001010001110001101" , -- ADDR 12
			"00000000000000000110100100101110" , -- ADDR 13
			"00000000000000001000110010101110" , -- ADDR 14
			"00000000000000000100100010101001" , -- ADDR 15
			"00000000000000000111011111010100" , -- ADDR 16
			"00000000000000000110101111000010" , -- ADDR 17
			"00000000000000001011001011100001" , -- ADDR 18
			"00000000000000000101000110010001" , -- ADDR 19
			"00000000000000000110100100101110" , -- ADDR 20
			"00000000000000000001101110011111" , -- ADDR 21
			"00000000000000000101010001010011" , -- ADDR 22
			"00000000000000000111000101001000" , -- ADDR 23
			"00000000000000001000000101010010" , -- ADDR 24
			"00000000000000000100100110110100" , -- ADDR 25
			"00000000000000000001111101111110" , -- ADDR 26
			"00000000000000000011111100011011" , -- ADDR 27
			"00000000000000000101001110000010" , -- ADDR 28
			"00000000000000000111111110001010" , -- ADDR 29
			"00000000000000000100001001101000" , -- ADDR 30
			"00000000000000000001011111000011" , -- ADDR 31
			"00000000000000001010011111001001" , -- ADDR 32
			"00000000000000000111011110010010" , -- ADDR 33
			"00000000000000000110101010110001" , -- ADDR 34
			"00000000000000000111100101011000" , -- ADDR 35
			"00000000000000000111011011001110" , -- ADDR 36
			"00000000000000000100100101100100" , -- ADDR 37
			"00000000000000001010100000100110" , -- ADDR 38
			"00000000000000001101101011100100" , -- ADDR 39
			"00000000000000001010110010101100" , -- ADDR 40
			"00000000000000001010111110010000" , -- ADDR 41
			"00000000000000001000010110000000" , -- ADDR 42
			"00000000000000001001001100011000" , -- ADDR 43
			"00000000000000001010010001000000" , -- ADDR 44
			"00000000000000000011011001101000" , -- ADDR 45
			"00000000000000000101101100011100" , -- ADDR 46
			"00000000000000000011000001010001" , -- ADDR 47
			"00000000000000000110011100100001" , -- ADDR 48
			"00000000000000000101111010001111" , -- ADDR 49
			"00000000000000000011011001000100" , -- ADDR 50
			"00000000000000000011101111000001" , -- ADDR 51
			"00000000000000001001000010010110" , -- ADDR 52
			"00000000000000000101001000100000" , -- ADDR 53
			"00000000000000000110110110100111" , -- ADDR 54
			"00000000000000001000100001110000" , -- ADDR 55
			"00000000000000000101011010111100" , -- ADDR 56
			"00000000000000000011111110010111" , -- ADDR 57
			"00000000000000000110110110100111" , -- ADDR 58
			"00000000000000000010100110000110" , -- ADDR 59
			"00000000000000000110000010110111" , -- ADDR 60
			"00000000000000001100001111001000" , -- ADDR 61
			"00000000000000001001001100011000" , -- ADDR 62
			"00000000000000001000101010001100" , -- ADDR 63
			"00000000000000000010000101100000" , -- ADDR 64
			"00000000000000001000010100001011" , -- ADDR 65
			"00000000000000001000101111000001" , -- ADDR 66
			"00000000000000001100011011100000" , -- ADDR 67
			"00000000000000000010111100001010" , -- ADDR 68
			"00000000000000000011100110101101" , -- ADDR 69
			"00000000000000000010100110000110" , -- ADDR 70
			"00000000000000001000010010100100" , -- ADDR 71
			"00000000000000001010000010010110" , -- ADDR 72
			"00000000000000001010100110011001" , -- ADDR 73
			"00000000000000000111000110001101" , -- ADDR 74
			"00000000000000000100101001010010" , -- ADDR 75
			"00000000000000000100101000011110" , -- ADDR 76
			"00000000000000000010001101011111" , -- ADDR 77
			"00000000000000000101110011011010" , -- ADDR 78
			"00000000000000000101101100011100" , -- ADDR 79
			"00000000000000000010110010001010" , -- ADDR 80
			"00000000000000001001100011001011" , -- ADDR 81
			"00000000000000000100111000100000" , -- ADDR 82
			"00000000000000000100101010100001" , -- ADDR 83
			"00000000000000000101111101011101" , -- ADDR 84
			"00000000000000000111110010100010" , -- ADDR 85
			"00000000000000000011100011100000" , -- ADDR 86
			"00000000000000001000101001110000" , -- ADDR 87
			"00000000000000001111000001010010" , -- ADDR 88
			"00000000000000001100010100010000" , -- ADDR 89
			"00000000000000001011101110001010" , -- ADDR 90
			"00000000000000001011010110010111" , -- ADDR 91
			"00000000000000001001100000100101" , -- ADDR 92
			"00000000000000001001110101000110" , -- ADDR 93
			"00000000000000000100110100001011" , -- ADDR 94
			"00000000000000000111001011100011" , -- ADDR 95
			"00000000000000000110000010100011" , -- ADDR 96
			"00000000000000000101001000100000" , -- ADDR 97
			"00000000000000000011011001000100" , -- ADDR 98
			"00000000000000000101001000100000" , -- ADDR 99
			"00000000000000001100001000001111" , -- ADDR 100
			"00000000000000001000110011011000" , -- ADDR 101
			"00000000000000001000101000011011" , -- ADDR 102
			"00000000000000001000100011000110" , -- ADDR 103
			"00000000000000000101001001100111" , -- ADDR 104
			"00000000000000000111100100011000" , -- ADDR 105
			"00000000000000001010100000000100" , -- ADDR 106
			"00000000000000000110000111111000" , -- ADDR 107
			"00000000000000001001010110000011" , -- ADDR 108
			"00000000000000001110111010010010" , -- ADDR 109
			"00000000000000001011001001010011" , -- ADDR 110
			"00000000000000001100010110100100" , -- ADDR 111
			"00000000000000000101100111011000" , -- ADDR 112
			"00000000000000001011101110010101" , -- ADDR 113
			"00000000000000001011011010100011" , -- ADDR 114
			"00000000000000001111101011001011" , -- ADDR 115
			"00000000000000000001111010000010" , -- ADDR 116
			"00000000000000000101111001100110" , -- ADDR 117
			"00000000000000000010111110101111" , -- ADDR 118
			"00000000000000001000111101000010" , -- ADDR 119
			"00000000000000001011001000100111" , -- ADDR 120
			"00000000000000001100101100000011" , -- ADDR 121
			"00000000000000000110001011100110" , -- ADDR 122
			"00000000000000000110101001000011" , -- ADDR 123
			"00000000000000000010010100001111" , -- ADDR 124
			"00000000000000000100001011000000" , -- ADDR 125
			"00000000000000001001001001101011" , -- ADDR 126
			"00000000000000000011110111000011" , -- ADDR 127
			"00000000000000000101100100010100" , -- ADDR 128
			"00000000000000001101010000111100" , -- ADDR 129
			"00000000000000000111111000011000" , -- ADDR 130
			"00000000000000000010011101000010" , -- ADDR 131
			"00000000000000000010111100110011" , -- ADDR 132
			"00000000000000001011010110110111" , -- ADDR 133
			"00000000000000000111010010001001" , -- ADDR 134
			"00000000000000001100000101011001" , -- ADDR 135
			"00000000000000010010001110011101" , -- ADDR 136
			"00000000000000001111011000111000" , -- ADDR 137
			"00000000000000001111001100111010" , -- ADDR 138
			"00000000000000001011011110011000" , -- ADDR 139
			"00000000000000001101000111010000" , -- ADDR 140
			"00000000000000001101100011110111" , -- ADDR 141
			"00000000000000000111110100010000" , -- ADDR 142
			"00000000000000001010001110001101" , -- ADDR 143
			"00000000000000000110111100101100" , -- ADDR 144
			"00000000000000001000110101111110" , -- ADDR 145
			"00000000000000000110101010011111" , -- ADDR 146
			"00000000000000000111111100101110" , -- ADDR 147
			"00000000000000000100111110101100" , -- ADDR 148
			"00000000000000000101001000100000" , -- ADDR 149
			"00000000000000001001000100000001" , -- ADDR 150
			"00000000000000001001001100001011" , -- ADDR 151
			"00000000000000000111111111110101" , -- ADDR 152
			"00000000000000000111101010101001" , -- ADDR 153
			"00000000000000000110100000000011" , -- ADDR 154
			"00000000000000000011000011110010" , -- ADDR 155
			"00000000000000000011101010111001" , -- ADDR 156
			"00000000000000000100010111100001" , -- ADDR 157
			"00000000000000000100100110110100" , -- ADDR 158
			"00000000000000001000101000001101" , -- ADDR 159
			"00000000000000000001110111000000" , -- ADDR 160
			"00000000000000000001110111000000" , -- ADDR 161
			"00000000000000000011100110101101" , -- ADDR 162
			"00000000000000001011111100010110" , -- ADDR 163
			"00000000000000001010111110010000" , -- ADDR 164
			"00000000000000001001010001111101" , -- ADDR 165
			"00000000000000000111101000011001" , -- ADDR 166
			"00000000000000000110111111011100" , -- ADDR 167
			"00000000000000000100010100011100" , -- ADDR 168
			"00000000000000001010011001010011" , -- ADDR 169
			"00000000000000000101111001100110" , -- ADDR 170
			"00000000000000001011011110100011" , -- ADDR 171
			"00000000000000001010101110000101" , -- ADDR 172
			"00000000000000001001010001111101" , -- ADDR 173
			"00000000000000001011010010011111" , -- ADDR 174
			"00000000000000000110100100011011" , -- ADDR 175
			"00000000000000000111011101000001" , -- ADDR 176
			"00000000000000001010001001111001" , -- ADDR 177
			"00000000000000001101101010100101" , -- ADDR 178
			"00000000000000001110110110001011" , -- ADDR 179
			"00000000000000000011000101101001" , -- ADDR 180
			"00000000000000000110011111001011" , -- ADDR 181
			"00000000000000001001111001001010" , -- ADDR 182
			"00000000000000000110000110101000" , -- ADDR 183
			"00000000000000000011010010001110" , -- ADDR 184
			"00000000000000000011111010011111" , -- ADDR 185
			"00000000000000001001111110010101" , -- ADDR 186
			"00000000000000000011101000010010" , -- ADDR 187
			"00000000000000000110000100000111" , -- ADDR 188
			"00000000000000000100010100011100" , -- ADDR 189
			"00000000000000000001111010000010" , -- ADDR 190
			"00000000000000000111001011110100" , -- ADDR 191
			"00000000000000000110110110100111" , -- ADDR 192
			"00000000000000001001001100001011" , -- ADDR 193
			"00000000000000000100001100110101" , -- ADDR 194
			"00000000000000000110001110010111" , -- ADDR 195
			"00000000000000001001110100100000" , -- ADDR 196
			"00000000000000001000000111011010" , -- ADDR 197
			"00000000000000000011000001010001" , -- ADDR 198
			"00000000000000000011011110000101" , -- ADDR 199
			"00000000000000000010101110101100" , -- ADDR 200
			"00000000000000000010010000000100" , -- ADDR 201
			"00000000000000001000101000011011" , -- ADDR 202
			"00000000000000000111011011111111" , -- ADDR 203
			"00000000000000000011100011100000" , -- ADDR 204
			"00000000000000000011111110010111" , -- ADDR 205
			"00000000000000000011100110101101" , -- ADDR 206
			"00000000000000000101101010011011" , -- ADDR 207
			"00000000000000000111110010100010" , -- ADDR 208
			"00000000000000000111111111110101" , -- ADDR 209
			"00000000000000000110000111100100" , -- ADDR 210
			"00000000000000000110100111000010" , -- ADDR 211
			"00000000000000001000110100011101" , -- ADDR 212
			"00000000000000001001011110110001" , -- ADDR 213
			"00000000000000001000010010100100" , -- ADDR 214
			"00000000000000001001110011100010" , -- ADDR 215
			"00000000000000000101000001101111" , -- ADDR 216
			"00000000000000001001000100000001" , -- ADDR 217
			"00000000000000000110001101110000" , -- ADDR 218
			"00000000000000000100011101001000" , -- ADDR 219
			"00000000000000001001100011001011" , -- ADDR 220
			"00000000000000000011111011111101" , -- ADDR 221
			"00000000000000000101000110010001" , -- ADDR 222
			"00000000000000000101001011011101" , -- ADDR 223
			"00000000000000001001101011101101" , -- ADDR 224
			"00000000000000001011000011011101" , -- ADDR 225
			"00000000000000000010110000110010" , -- ADDR 226
			"00000000000000000001101110011111" , -- ADDR 227
			"00000000000000000101111010001111" , -- ADDR 228
			"00000000000000001010010111000110" , -- ADDR 229
			"00000000000000000111111110111000" , -- ADDR 230
			"00000000000000000110101111000010" , -- ADDR 231
			"00000000000000001011111010011011" , -- ADDR 232
			"00000000000000000100011001101100" , -- ADDR 233
			"00000000000000000100111000111001" , -- ADDR 234
			"00000000000000000010111100001010" , -- ADDR 235
			"00000000000000000011101100011101" , -- ADDR 236
			"00000000000000000111000111100011" , -- ADDR 237
			"00000000000000000010000000110110" , -- ADDR 238
			"00000000000000000100010000111000" , -- ADDR 239
			"00000000000000000011011100111110" , -- ADDR 240
			"00000000000000000100000001101100" , -- ADDR 241
			"00000000000000000100011001101100" , -- ADDR 242
			"00000000000000001000010011011111" , -- ADDR 243
			"00000000000000001001101100010011" , -- ADDR 244
			"00000000000000000101010101010000" , -- ADDR 245
			"00000000000000000100011001101100" , -- ADDR 246
			"00000000000000000110101001000011" , -- ADDR 247
			"00000000000000000010100000111000" , -- ADDR 248
			"00000000000000001000011010000110" , -- ADDR 249
			"00000000000000000111101101010111" , -- ADDR 250
			"00000000000000000110000010100011" , -- ADDR 251
			"00000000000000000011100011100000" , -- ADDR 252
			"00000000000000001000100001110000" , -- ADDR 253
			"00000000000000001001001100001011" , -- ADDR 254
			"00000000000000001010000101011000" , -- ADDR 255
			"00000000000000000101101011011011" , -- ADDR 256
			"00000000000000000010101110101100" , -- ADDR 257
			"00000000000000000011011001101000" , -- ADDR 258
			"00000000000000000100000100000011" , -- ADDR 259
			"00000000000000000101010101010000" , -- ADDR 260
			"00000000000000000010001101011111" , -- ADDR 261
			"00000000000000000111010000100100" , -- ADDR 262
			"00000000000000001001000010010110" , -- ADDR 263
			"00000000000000001010010001001011" , -- ADDR 264
			"00000000000000000110101001000011" , -- ADDR 265
			"00000000000000000100001010000101" , -- ADDR 266
			"00000000000000001010111001101110" , -- ADDR 267
			"00000000000000001010010110001011" , -- ADDR 268
			"00000000000000001010101111101011" , -- ADDR 269
			"00000000000000001011100100110101" , -- ADDR 270
			"00000000000000000110101010110001" , -- ADDR 271
			"00000000000000000110100011010001" , -- ADDR 272
			"00000000000000001100001000001111" , -- ADDR 273
			"00000000000000001010101111101011" , -- ADDR 274
			"00000000000000000111110011010001" , -- ADDR 275
			"00000000000000001001000010001000" , -- ADDR 276
			"00000000000000000101101100110001" , -- ADDR 277
			"00000000000000001000000111011010" , -- ADDR 278
			"00000000000000001010000010111010" , -- ADDR 279
			"00000000000000000011010100100001" , -- ADDR 280
			"00000000000000000011110010100100" , -- ADDR 281
			"00000000000000000010001011110000" , -- ADDR 282
			"00000000000000001000000011110111" , -- ADDR 283
			"00000000000000001000111000110001" , -- ADDR 284
			"00000000000000000010110010001010" , -- ADDR 285
			"00000000000000000011011011010100" , -- ADDR 286
			"00000000000000001011010000010010" , -- ADDR 287
			"00000000000000001101001100010101" , -- ADDR 288
			"00000000000000001000001000010110" , -- ADDR 289
			"00000000000000001000010011011111" , -- ADDR 290
			"00000000000000001001101110101010" , -- ADDR 291
			"00000000000000000101010001010011" , -- ADDR 292
			"00000000000000001100011000000111" , -- ADDR 293
			"00000000000000001010000101111100" , -- ADDR 294
			"00000000000000001010000100001111" , -- ADDR 295
			"00000000000000000111010100110000" , -- ADDR 296
			"00000000000000001100001111110000" , -- ADDR 297
			"00000000000000001001110101110111" , -- ADDR 298
			"00000000000000001100000111111011" , -- ADDR 299
			"00000000000000000110010001101110" , -- ADDR 300
			"00000000000000000001011111000011" , -- ADDR 301
			"00000000000000000011011110000101" , -- ADDR 302
			"00000000000000000110100100101110" , -- ADDR 303
			"00000000000000000010101110101100" , -- ADDR 304
			"00000000000000000100110110001001" , -- ADDR 305
			"00000000000000000110011011000010" , -- ADDR 306
			"00000000000000001010101010001010" , -- ADDR 307
			"00000000000000001101010100100010" , -- ADDR 308
			"00000000000000000101000110010001" , -- ADDR 309
			"00000000000000000110100110001011" , -- ADDR 310
			"00000000000000001110101111111111" , -- ADDR 311
			"00000000000000001101000000000110" , -- ADDR 312
			"00000000000000001010111111001000" , -- ADDR 313
			"00000000000000001011010100110110" , -- ADDR 314
			"00000000000000001010101010001010" , -- ADDR 315
			"00000000000000001001101010101110" , -- ADDR 316
			"00000000000000001111100100100101" , -- ADDR 317
			"00000000000000001110001110001001" , -- ADDR 318
			"00000000000000001011010111000010" , -- ADDR 319
			"00000000000000001100111110011111" , -- ADDR 320
			"00000000000000000010111100001010" , -- ADDR 321
			"00000000000000001100001001000001" , -- ADDR 322
			"00000000000000001110000000101001" , -- ADDR 323
			"00000000000000000110111010001110" , -- ADDR 324
			"00000000000000000111110100010000" , -- ADDR 325
			"00000000000000000010110000110010" , -- ADDR 326
			"00000000000000001011011010100011" , -- ADDR 327
			"00000000000000001011011100011000" , -- ADDR 328
			"00000000000000000110011100110100" , -- ADDR 329
			"00000000000000001000101111011101" , -- ADDR 330
			"00000000000000001011001000110010" , -- ADDR 331
			"00000000000000000101110010011011" , -- ADDR 332
			"00000000000000000111010100110000" , -- ADDR 333
			"00000000000000001011000010100110" , -- ADDR 334
			"00000000000000000110101111000010" , -- ADDR 335
			"00000000000000001011010010111111" , -- ADDR 336
			"00000000000000000111010000000010" , -- ADDR 337
			"00000000000000001001100100100101" , -- ADDR 338
			"00000000000000000111110111001010" , -- ADDR 339
			"00000000000000001100101111101010" , -- ADDR 340
			"00000000000000000110011011000010" , -- ADDR 341
			"00000000000000001001000000011100" , -- ADDR 342
			"00000000000000000010111100110011" , -- ADDR 343
			"00000000000000000011110111000011" , -- ADDR 344
			"00000000000000000110000111111000" , -- ADDR 345
			"00000000000000001000010010010101" , -- ADDR 346
			"00000000000000000001110000101011" , -- ADDR 347
			"00000000000000000011011011010100" , -- ADDR 348
			"00000000000000000011001011001000" , -- ADDR 349
			"00000000000000000111011011001110" , -- ADDR 350
			"00000000000000001010110010101100" , -- ADDR 351
			"00000000000000000010010000000100" , -- ADDR 352
			"00000000000000000100010000111000" , -- ADDR 353
			"00000000000000001101001101101000" , -- ADDR 354
			"00000000000000001010001011111101" , -- ADDR 355
			"00000000000000000111100100101000" , -- ADDR 356
			"00000000000000000111111111110101" , -- ADDR 357
			"00000000000000001001110001001100" , -- ADDR 358
			"00000000000000000111011011001110" , -- ADDR 359
			"00000000000000001101010110110100" , -- ADDR 360
			"00000000000000001111000100101101" , -- ADDR 361
			"00000000000000001100000111111011" , -- ADDR 362
			"00000000000000001100111011011001" , -- ADDR 363
			"00000000000000000110010111011101" , -- ADDR 364
			"00000000000000001011011110100011" , -- ADDR 365
			"00000000000000001100110110000100" , -- ADDR 366
			"00000000000000000101100111101110" , -- ADDR 367
			"00000000000000000111011110000010" , -- ADDR 368
			"00000000000000000010010000000100" , -- ADDR 369
			"00000000000000001001010001111101" , -- ADDR 370
			"00000000000000001000101000011011" , -- ADDR 371
			"00000000000000000101011000000111" , -- ADDR 372
			"00000000000000000010111100001010" , -- ADDR 373
			"00000000000000000011001000000110" , -- ADDR 374
			"00000000000000000101001000100000" , -- ADDR 375
			"00000000000000001011101000111100" , -- ADDR 376
			"00000000000000001010000000101000" , -- ADDR 377
			"00000000000000000101101100110001" , -- ADDR 378
			"00000000000000000001111101000000" , -- ADDR 379
			"00000000000000000110100100101110" , -- ADDR 380
			"00000000000000001000100010111000" , -- ADDR 381
			"00000000000000001010101100110101" , -- ADDR 382
			"00000000000000000110001110010111" , -- ADDR 383
			"00000000000000000011010010001110" , -- ADDR 384
			"00000000000000000110010110010000" , -- ADDR 385
			"00000000000000001010100100000011" , -- ADDR 386
			"00000000000000001011101100110111" , -- ADDR 387
			"00000000000000001011000011011101" , -- ADDR 388
			"00000000000000001010100000000100" , -- ADDR 389
			"00000000000000000110100000000011" , -- ADDR 390
			"00000000000000001000100101100011" , -- ADDR 391
			"00000000000000000011111100011011" , -- ADDR 392
			"00000000000000000010000100100101" , -- ADDR 393
			"00000000000000001001100001011000" , -- ADDR 394
			"00000000000000000100101010100001" , -- ADDR 395
			"00000000000000000101110011011010" , -- ADDR 396
			"00000000000000000010001100101000" , -- ADDR 397
			"00000000000000000111101110000111" , -- ADDR 398
			"00000000000000001001001100001011" , -- ADDR 399
			"00000000000000000101100100101001" , -- ADDR 400
			"00000000000000000001110001110000" , -- ADDR 401
			"00000000000000000100101101110001" , -- ADDR 402
			"00000000000000001101001110111011" , -- ADDR 403
			"00000000000000001010111110010000" , -- ADDR 404
			"00000000000000001001011011001001" , -- ADDR 405
			"00000000000000001101101111101111" , -- ADDR 406
			"00000000000000000110111100001001" , -- ADDR 407
			"00000000000000000110011100110100" , -- ADDR 408
			"00000000000000000101000110010001" , -- ADDR 409
			"00000000000000000110100110001011" , -- ADDR 410
			"00000000000000001000100000001100" , -- ADDR 411
			"00000000000000000001100100000011" , -- ADDR 412
			"00000000000000000001011000011001" , -- ADDR 413
			"00000000000000000101101000101111" , -- ADDR 414
			"00000000000000000101010110101100" , -- ADDR 415
			"00000000000000000101100100101001" , -- ADDR 416
			"00000000000000001011010001011110" , -- ADDR 417
			"00000000000000001010110100000110" , -- ADDR 418
			"00000000000000000011110111000011" , -- ADDR 419
			"00000000000000000100111000111001" , -- ADDR 420
			"00000000000000000101111000010011" , -- ADDR 421
			"00000000000000001000110011011000" , -- ADDR 422
			"00000000000000001001011110110001" , -- ADDR 423
			"00000000000000001001001001101011" , -- ADDR 424
			"00000000000000000101110010011011" , -- ADDR 425
			"00000000000000001001000011110100" , -- ADDR 426
			"00000000000000001100010000100010" , -- ADDR 427
			"00000000000000001100111100010001" , -- ADDR 428
			"00000000000000001011100001000010" , -- ADDR 429
			"00000000000000001100111000100101" , -- ADDR 430
			"00000000000000001000010110011101" , -- ADDR 431
			"00000000000000001011011001100010" , -- ADDR 432
			"00000000000000000110110011110101" , -- ADDR 433
			"00000000000000000010010000000100" , -- ADDR 434
			"00000000000000001100001101010000" , -- ADDR 435
			"00000000000000000110111000010010" , -- ADDR 436
			"00000000000000000010111100110011" , -- ADDR 437
			"00000000000000000011110100000100" , -- ADDR 438
			"00000000000000001010100110011001" , -- ADDR 439
			"00000000000000001100000101000101" , -- ADDR 440
			"00000000000000000100101001010010" , -- ADDR 441
			"00000000000000000011101110000000" , -- ADDR 442
			"00000000000000000010011100010000" , -- ADDR 443
			"00000000000000001011110100000000" , -- ADDR 444
			"00000000000000001010000011101011" , -- ADDR 445
			"00000000000000000111110011010001" , -- ADDR 446
			"00000000000000001111010111111000" , -- ADDR 447
			"00000000000000000101010101010000" , -- ADDR 448
			"00000000000000000011111110010111" , -- ADDR 449
			"00000000000000000110011000111101" , -- ADDR 450
			"00000000000000000110111001000111" , -- ADDR 451
			"00000000000000001010011100110010" , -- ADDR 452
			"00000000000000000001110111000000" , -- ADDR 453
			"00000000000000000100000101111011" , -- ADDR 454
			"00000000000000000110111010100000" , -- ADDR 455
			"00000000000000000011011110000101" , -- ADDR 456
			"00000000000000001001110101110111" , -- ADDR 457
			"00000000000000000111010101000001" , -- ADDR 458
			"00000000000000000110010001101110" , -- ADDR 459
			"00000000000000000010011100010000" , -- ADDR 460
			"00000000000000000101101110000111" , -- ADDR 461
			"00000000000000000110011010001001" , -- ADDR 462
			"00000000000000001001110101110111" , -- ADDR 463
			"00000000000000000101100010010000" , -- ADDR 464
			"00000000000000000100111000111001" , -- ADDR 465
			"00000000000000000011111010000000" , -- ADDR 466
			"00000000000000000111011101000001" , -- ADDR 467
			"00000000000000001000101110010111" , -- ADDR 468
			"00000000000000001000100100111000" , -- ADDR 469
			"00000000000000000111100010100111" , -- ADDR 470
			"00000000000000000011011001000100" , -- ADDR 471
			"00000000000000000110010110100011" , -- ADDR 472
			"00000000000000000100010000111000" , -- ADDR 473
			"00000000000000000101001100001100" , -- ADDR 474
			"00000000000000000110111100011011" , -- ADDR 475
			"00000000000000000001100100000011" , -- ADDR 476
			"00000000000000000111101000011001" , -- ADDR 477
			"00000000000000000101000010001000" , -- ADDR 478
			"00000000000000000111010000100100" , -- ADDR 479
			"00000000000000001000100010111000" , -- ADDR 480
			"00000000000000000101001111011111" , -- ADDR 481
			"00000000000000000001101000110100" , -- ADDR 482
			"00000000000000000111100101011000" , -- ADDR 483
			"00000000000000001100011011110011" , -- ADDR 484
			"00000000000000001001110001000000" , -- ADDR 485
			"00000000000000001001001001000011" , -- ADDR 486
			"00000000000000001010101000101110" , -- ADDR 487
			"00000000000000000110111111011100" , -- ADDR 488
			"00000000000000000111100110101001" , -- ADDR 489
			"00000000000000000010011111010110" , -- ADDR 490
			"00000000000000000100101100100011" , -- ADDR 491
			"00000000000000000101011000000111" , -- ADDR 492
			"00000000000000000011011111101110" , -- ADDR 493
			"00000000000000000011100011100000" , -- ADDR 494
			"00000000000000000010111100001010" , -- ADDR 495
			"00000000000000000110100100101110" , -- ADDR 496
			"00000000000000000101001111011111" , -- ADDR 497
			"00000000000000000100000101111011" , -- ADDR 498
			"00000000000000000101100100111111" , -- ADDR 499
			"00000000000000000010011001111001" , -- ADDR 500
			"00000000000000000011011011010100" , -- ADDR 501
			"00000000000000000110011000111101" , -- ADDR 502
			"00000000000000001000111110100010" , -- ADDR 503
			"00000000000000000111111100111101" , -- ADDR 504
			"00000000000000000110101010110001" , -- ADDR 505
			"00000000000000000111000111100011" , -- ADDR 506
			"00000000000000000111011100010000" , -- ADDR 507
			"00000000000000000110000010100011" , -- ADDR 508
			"00000000000000001000110101111110" , -- ADDR 509
			"00000000000000000011111010011111" , -- ADDR 510
			"00000000000000001001000010001000" , -- ADDR 511
			"00000000000000000111101010011001" , -- ADDR 512
			"00000000000000000110101101000011" , -- ADDR 513
			"00000000000000001001001001101011" , -- ADDR 514
			"00000000000000000011110100100100" , -- ADDR 515
			"00000000000000000110100000000011" , -- ADDR 516
			"00000000000000000111010101000001" , -- ADDR 517
			"00000000000000001010101101000001" , -- ADDR 518
			"00000000000000001011111100010110" , -- ADDR 519
			"00000000000000000010011101000010" , -- ADDR 520
			"00000000000000000011011111101110" , -- ADDR 521
			"00000000000000000111111111110101" , -- ADDR 522
			"00000000000000001000111110100010" , -- ADDR 523
			"00000000000000000110010011001111" , -- ADDR 524
			"00000000000000000101111001100110" , -- ADDR 525
			"00000000000000001010000100001111" , -- ADDR 526
			"00000000000000000100001010000101" , -- ADDR 527
			"00000000000000000101101101110001" , -- ADDR 528
			"00000000000000000001101110011111" , -- ADDR 529
			"00000000000000000001011101110000" , -- ADDR 530
			"00000000000000000101110011011010" , -- ADDR 531
			"00000000000000000100010000111000" , -- ADDR 532
			"00000000000000000110001110010111" , -- ADDR 533
			"00000000000000000001111101111110" , -- ADDR 534
			"00000000000000000100011111010001" , -- ADDR 535
			"00000000000000000111111000011000" , -- ADDR 536
			"00000000000000001100000111110001" , -- ADDR 537
			"00000000000000000101011001001011" , -- ADDR 538
			"00000000000000000011100001010110" , -- ADDR 539
			"00000000000000000011100001010110" , -- ADDR 540
			"00000000000000001111000010010011" , -- ADDR 541
			"00000000000000001110100001011001" , -- ADDR 542
			"00000000000000001011111100010110" , -- ADDR 543
			"00000000000000001000010000101110" , -- ADDR 544
			"00000000000000000110101000011110" , -- ADDR 545
			"00000000000000000011001101100001" , -- ADDR 546
			"00000000000000001011110010101101" , -- ADDR 547
			"00000000000000001000010010110011" , -- ADDR 548
			"00000000000000001101110100111111" , -- ADDR 549
			"00000000000000001110000110101111" , -- ADDR 550
			"00000000000000001100111100101110" , -- ADDR 551
			"00000000000000001101010010000110" , -- ADDR 552
			"00000000000000001001100011001011" , -- ADDR 553
			"00000000000000001010101010001010" , -- ADDR 554
			"00000000000000001101110011111001" , -- ADDR 555
			"00000000000000010000101110011001" , -- ADDR 556
			"00000000000000010001110001100001" , -- ADDR 557
			"00000000000000000110101000011110" , -- ADDR 558
			"00000000000000001010000100001111" , -- ADDR 559
			"00000000000000001101011010000110" , -- ADDR 560
			"00000000000000000100101000111000" , -- ADDR 561
			"00000000000000000010010011011010" , -- ADDR 562
			"00000000000000000101010110101100" , -- ADDR 563
			"00000000000000001001100001011000" , -- ADDR 564
			"00000000000000000110100100101110" , -- ADDR 565
			"00000000000000001001000100101010" , -- ADDR 566
			"00000000000000000111011011001110" , -- ADDR 567
			"00000000000000000101001011000110" , -- ADDR 568
			"00000000000000001000110011011000" , -- ADDR 569
			"00000000000000001010100001100001" , -- ADDR 570
			"00000000000000001100110010101001" , -- ADDR 571
			"00000000000000000111000111100011" , -- ADDR 572
			"00000000000000001000101000111000" , -- ADDR 573
			"00000000000000001001110001001100" , -- ADDR 574
			"00000000000000000101111010001111" , -- ADDR 575
			"00000000000000000010100000111000" , -- ADDR 576
			"00000000000000000111000101011001" , -- ADDR 577
			"00000000000000001011101010010000" , -- ADDR 578
			"00000000000000001100001101010000" , -- ADDR 579
			"00000000000000001000001100000101" , -- ADDR 580
			"00000000000000000011110010100100" , -- ADDR 581
			"00000000000000000010101000010010" , -- ADDR 582
			"00000000000000000001100100000011" , -- ADDR 583
			"00000000000000000111010101000001" , -- ADDR 584
			"00000000000000000100101000011110" , -- ADDR 585
			"00000000000000001001101110010001" , -- ADDR 586
			"00000000000000001011010100110110" , -- ADDR 587
			"00000000000000001011110100000000" , -- ADDR 588
			"00000000000000001000111110111101" , -- ADDR 589
			"00000000000000000110011011000010" , -- ADDR 590
			"00000000000000001011011001100010" , -- ADDR 591
			"00000000000000001100001010011100" , -- ADDR 592
			"00000000000000001101001111010111" , -- ADDR 593
			"00000000000000001110000101101010" , -- ADDR 594
			"00000000000000000110111001111100" , -- ADDR 595
			"00000000000000001000001111000110" , -- ADDR 596
			"00000000000000001101001110111011" , -- ADDR 597
			"00000000000000001000111101000010" , -- ADDR 598
			"00000000000000000110000111111000" , -- ADDR 599
			"00000000000000001000000111011010" , -- ADDR 600
			"00000000000000000101101000101111" , -- ADDR 601
			"00000000000000000111111011000010" , -- ADDR 602
			"00000000000000001010001110001101" , -- ADDR 603
			"00000000000000000100111100000000" , -- ADDR 604
			"00000000000000000100000000010001" , -- ADDR 605
			"00000000000000000100011111010001" , -- ADDR 606
			"00000000000000001001011011100010" , -- ADDR 607
			"00000000000000001010110011111011" , -- ADDR 608
			"00000000000000000100011010111111" , -- ADDR 609
			"00000000000000000111001111110010" , -- ADDR 610
			"00000000000000000010110010001010" , -- ADDR 611
			"00000000000000000110001110010111" , -- ADDR 612
			"00000000000000000101101010011011" , -- ADDR 613
			"00000000000000001011011101101101" , -- ADDR 614
			"00000000000000001000111110100010" , -- ADDR 615
			"00000000000000001010000111011101" , -- ADDR 616
			"00000000000000001011001000110010" , -- ADDR 617
			"00000000000000001011001000100111" , -- ADDR 618
			"00000000000000001000111000110001" , -- ADDR 619
			"00000000000000001100111000100101" , -- ADDR 620
			"00000000000000000111111100101110" , -- ADDR 621
			"00000000000000001100100100010110" , -- ADDR 622
			"00000000000000001001011110110001" , -- ADDR 623
			"00000000000000000110000000010101" , -- ADDR 624
			"00000000000000001100111100010001" , -- ADDR 625
			"00000000000000000111010101110011" , -- ADDR 626
			"00000000000000000010110110001110" , -- ADDR 627
			"00000000000000000111011000011000" , -- ADDR 628
			"00000000000000001101000111010000" , -- ADDR 629
			"00000000000000001110100001011001" , -- ADDR 630
			"00000000000000000001110000101011" , -- ADDR 631
			"00000000000000000101001000100000" , -- ADDR 632
			"00000000000000000101100111101110" , -- ADDR 633
			"00000000000000000111111100111101" , -- ADDR 634
			"00000000000000000110010110100011" , -- ADDR 635
			"00000000000000000011111100011011" , -- ADDR 636
			"00000000000000001101111100110100" , -- ADDR 637
			"00000000000000000001011111000011" , -- ADDR 638
			"00000000000000000001101000110100" , -- ADDR 639
			"00000000000000000101101100110001" , -- ADDR 640
			"00000000000000000100101111011000" , -- ADDR 641
			"00000000000000001001111001001010" , -- ADDR 642
			"00000000000000000100001001001011" , -- ADDR 643
			"00000000000000000111000101001000" , -- ADDR 644
			"00000000000000000110000010100011" , -- ADDR 645
			"00000000000000000111100001010110" , -- ADDR 646
			"00000000000000001000110000111111" , -- ADDR 647
			"00000000000000001011101110001010" , -- ADDR 648
			"00000000000000000100010100111000" , -- ADDR 649
			"00000000000000000010011101000010" , -- ADDR 650
			"00000000000000000100100110110100" , -- ADDR 651
			"00000000000000001001100111100011" , -- ADDR 652
			"00000000000000001011000100101010" , -- ADDR 653
			"00000000000000001011000000101100" , -- ADDR 654
			"00000000000000001000111110111101" , -- ADDR 655
			"00000000000000000101101000101111" , -- ADDR 656
			"00000000000000000110101101111010" , -- ADDR 657
			"00000000000000000010010000000100" , -- ADDR 658
			"00000000000000000011101110000000" , -- ADDR 659
			"00000000000000000111110000010101" , -- ADDR 660
			"00000000000000000011101000010010" , -- ADDR 661
			"00000000000000000111101101010111" , -- ADDR 662
			"00000000000000000010111100001010" , -- ADDR 663
			"00000000000000000101111001100110" , -- ADDR 664
			"00000000000000000111010110000011" , -- ADDR 665
			"00000000000000000110101111000010" , -- ADDR 666
			"00000000000000000010010000000100" , -- ADDR 667
			"00000000000000000110100100101110" , -- ADDR 668
			"00000000000000001110010011101000" , -- ADDR 669
			"00000000000000001011110011110110" , -- ADDR 670
			"00000000000000001010101101000001" , -- ADDR 671
			"00000000000000001100110001100110" , -- ADDR 672
			"00000000000000001000010100001011" , -- ADDR 673
			"00000000000000001000001101001111" , -- ADDR 674
			"00000000000000000100111010000100" , -- ADDR 675
			"00000000000000000110111100101100" , -- ADDR 676
			"00000000000000000111011011001110" , -- ADDR 677
			"00000000000000000011010100100001" , -- ADDR 678
			"00000000000000000001011000011001" , -- ADDR 679
			"00000000000000000101011000000111" , -- ADDR 680
			"00000000000000000011011100111110" , -- ADDR 681
			"00000000000000000100001100110101" , -- ADDR 682
			"00000000000000001011010000010010" , -- ADDR 683
			"00000000000000001001101110010001" , -- ADDR 684
			"00000000000000001001000100101010" , -- ADDR 685
			"00000000000000001000101110010111" , -- ADDR 686
			"00000000000000001000011101101110" , -- ADDR 687
			"00000000000000000110000110101000" , -- ADDR 688
			"00000000000000001010111111001000" , -- ADDR 689
			"00000000000000000110001001011011" , -- ADDR 690
			"00000000000000001011011011100011" , -- ADDR 691
			"00000000000000001001101110010001" , -- ADDR 692
			"00000000000000000111101000011001" , -- ADDR 693
			"00000000000000001011011111100010" , -- ADDR 694
			"00000000000000000110001110010111" , -- ADDR 695
			"00000000000000000101100111101110" , -- ADDR 696
			"00000000000000001000101001110000" , -- ADDR 697
			"00000000000000001100111110011111" , -- ADDR 698
			"00000000000000001110010000101100" , -- ADDR 699
			"00000000000000000001001111101011" , -- ADDR 700
			"00000000000000000101010010000001" , -- ADDR 701
			"00000000000000001000000011011001" , -- ADDR 702
			"00000000000000000110110010011011" , -- ADDR 703
			"00000000000000000100011001101100" , -- ADDR 704
			"00000000000000000011011111101110" , -- ADDR 705
			"00000000000000001011010111000010" , -- ADDR 706
			"00000000000000000010000101100000" , -- ADDR 707
			"00000000000000000100010100011100" , -- ADDR 708
			"00000000000000000100000101111011" , -- ADDR 709
			"00000000000000000010010000000100" , -- ADDR 710
			"00000000000000000111110100111110" , -- ADDR 711
			"00000000000000000101010001010011" , -- ADDR 712
			"00000000000000000111110111001010" , -- ADDR 713
			"00000000000000000100001101101111" , -- ADDR 714
			"00000000000000000100111110101100" , -- ADDR 715
			"00000000000000001011100001000010" , -- ADDR 716
			"00000000000000001011001101000011" , -- ADDR 717
			"00000000000000001000011101011111" , -- ADDR 718
			"00000000000000000101110111010101" , -- ADDR 719
			"00000000000000000101001000100000" , -- ADDR 720
			"00000000000000000010101110101100" , -- ADDR 721
			"00000000000000001000111000110001" , -- ADDR 722
			"00000000000000000100110110001001" , -- ADDR 723
			"00000000000000001010011100110010" , -- ADDR 724
			"00000000000000001010101010001010" , -- ADDR 725
			"00000000000000001010000111011101" , -- ADDR 726
			"00000000000000001010000011011111" , -- ADDR 727
			"00000000000000000110000001111010" , -- ADDR 728
			"00000000000000001001000010010110" , -- ADDR 729
			"00000000000000001010101111100000" , -- ADDR 730
			"00000000000000001101001101000011" , -- ADDR 731
			"00000000000000001110010000101100" , -- ADDR 732
			"00000000000000000100100010101001" , -- ADDR 733
			"00000000000000000110110110100111" , -- ADDR 734
			"00000000000000001011001001111111" , -- ADDR 735
			"00000000000000000111001101101011" , -- ADDR 736
			"00000000000000000100010000111000" , -- ADDR 737
			"00000000000000000101101100110001" , -- ADDR 738
			"00000000000000001000000111011010" , -- ADDR 739
			"00000000000000000101011010111100" , -- ADDR 740
			"00000000000000000111110001010100" , -- ADDR 741
			"00000000000000000011111100011011" , -- ADDR 742
			"00000000000000000001111101111110" , -- ADDR 743
			"00000000000000000101101101110001" , -- ADDR 744
			"00000000000000000111101010101001" , -- ADDR 745
			"00000000000000001001100100100101" , -- ADDR 746
			"00000000000000000011100110101101" , -- ADDR 747
			"00000000000000001111010111011000" , -- ADDR 748
			"00000000000000001101111001101011" , -- ADDR 749
			"00000000000000001100110111011001" , -- ADDR 750
			"00000000000000001010110001000110" , -- ADDR 751
			"00000000000000001001100110010111" , -- ADDR 752
			"00000000000000000110010001101110" , -- ADDR 753
			"00000000000000001101110110110010" , -- ADDR 754
			"00000000000000001001011111111110" , -- ADDR 755
			"00000000000000001111000101001110" , -- ADDR 756
			"00000000000000001101111010110001" , -- ADDR 757
			"00000000000000001011100000010111" , -- ADDR 758
			"00000000000000001110110111111110" , -- ADDR 759
			"00000000000000001010000110111000" , -- ADDR 760
			"00000000000000001000000101110000" , -- ADDR 761
			"00000000000000001100101100100000" , -- ADDR 762
			"00000000000000010001000101110111" , -- ADDR 763
			"00000000000000010010010101000001" , -- ADDR 764
			"00000000000000000101001000100000" , -- ADDR 765
			"00000000000000001001011110110001" , -- ADDR 766
			"00000000000000001011001111011011" , -- ADDR 767
			"00000000000000000010100110000110" , -- ADDR 768
			"00000000000000000001001110001000" , -- ADDR 769
			"00000000000000000010000101100000" , -- ADDR 770
			"00000000000000001100100110101000" , -- ADDR 771
			"00000000000000000100001011011101" , -- ADDR 772
			"00000000000000000110011000111101" , -- ADDR 773
			"00000000000000000111110111001010" , -- ADDR 774
			"00000000000000000101011111001000" , -- ADDR 775
			"00000000000000001010101010100001" , -- ADDR 776
			"00000000000000001001010010111111" , -- ADDR 777
			"00000000000000001100000001011100" , -- ADDR 778
			"00000000000000000111110010100010" , -- ADDR 779
			"00000000000000000100000101111011" , -- ADDR 780
			"00000000000000000011101010111001" , -- ADDR 781
			"00000000000000001010000000110100" , -- ADDR 782
			"00000000000000001100000011010110" , -- ADDR 783
			"00000000000000001101001001011100" , -- ADDR 784
			"00000000000000000111101110000111" , -- ADDR 785
			"00000000000000000111000001111000" , -- ADDR 786
			"00000000000000000100000100000011" , -- ADDR 787
			"00000000000000000010011101000010" , -- ADDR 788
			"00000000000000000111100100101000" , -- ADDR 789
			"00000000000000000101100100101001" , -- ADDR 790
			"00000000000000000101011111001000" , -- ADDR 791
			"00000000000000001100000001011100" , -- ADDR 792
			"00000000000000000110001011100110" , -- ADDR 793
			"00000000000000000001101110011111" , -- ADDR 794
			"00000000000000000011000011110010" , -- ADDR 795
			"00000000000000001010101100110101" , -- ADDR 796
			"00000000000000000110010101010110" , -- ADDR 797
			"00000000000000001010100000100110" , -- ADDR 798
			"00000000000000010001111101000011" , -- ADDR 799
			"00000000000000001111001110100010" , -- ADDR 800
			"00000000000000001110101001100000" , -- ADDR 801
			"00000000000000001100110001111001" , -- ADDR 802
			"00000000000000001100011001010110" , -- ADDR 803
			"00000000000000001100100001000000" , -- ADDR 804
			"00000000000000000111101010101001" , -- ADDR 805
			"00000000000000001010000100001111" , -- ADDR 806
			"00000000000000000111110110001100" , -- ADDR 807
			"00000000000000000111101001011001" , -- ADDR 808
			"00000000000000000101001000100000" , -- ADDR 809
			"00000000000000000111111011000010" , -- ADDR 810
			"00000000000000000110000110101000" , -- ADDR 811
			"00000000000000001011110100000000" , -- ADDR 812
			"00000000000000001101011010000110" , -- ADDR 813
			"00000000000000001101011101101001" , -- ADDR 814
			"00000000000000001010101001010000" , -- ADDR 815
			"00000000000000000111111100101110" , -- ADDR 816
			"00000000000000000111101010101001" , -- ADDR 817
			"00000000000000000001110000101011" , -- ADDR 818
			"00000000000000000011110010100100" , -- ADDR 819
			"00000000000000001000111110111101" , -- ADDR 820
			"00000000000000000101111100001011" , -- ADDR 821
			"00000000000000001000101111000001" , -- ADDR 822
			"00000000000000000010001101011111" , -- ADDR 823
			"00000000000000000101001000001000" , -- ADDR 824
			"00000000000000000110100110001011" , -- ADDR 825
			"00000000000000001000110011011000" , -- ADDR 826
			"00000000000000000100011111010001" , -- ADDR 827
			"00000000000000000110101000011110" , -- ADDR 828
			"00000000000000010000011101011001" , -- ADDR 829
			"00000000000000001110000101100001" , -- ADDR 830
			"00000000000000001100101100101010" , -- ADDR 831
			"00000000000000001110111010101010" , -- ADDR 832
			"00000000000000001010001110001101" , -- ADDR 833
			"00000000000000001001100111110000" , -- ADDR 834
			"00000000000000000111010111000110" , -- ADDR 835
			"00000000000000001001010110111000" , -- ADDR 836
			"00000000000000001001100100110001" , -- ADDR 837
			"00000000000000000100110101010111" , -- ADDR 838
			"00000000000000000001111010000010" , -- ADDR 839
			"00000000000000000111110100111110" , -- ADDR 840
			"00000000000000000110010110010000" , -- ADDR 841
			"00000000000000001000011000111110" , -- ADDR 842
			"00000000000000001001101110010001" , -- ADDR 843
			"00000000000000000100100010101001" , -- ADDR 844
			"00000000000000000011101010011000" , -- ADDR 845
			"00000000000000000010011101000010" , -- ADDR 846
			"00000000000000000100011110110110" , -- ADDR 847
			"00000000000000001000010011010000" , -- ADDR 848
			"00000000000000000011001011001000" , -- ADDR 849
			"00000000000000000010110110111001" , -- ADDR 850
			"00000000000000001011100001000010" , -- ADDR 851
			"00000000000000000111011110010010" , -- ADDR 852
			"00000000000000000101000110010001" , -- ADDR 853
			"00000000000000000101111001111011" , -- ADDR 854
			"00000000000000001000111000110001" , -- ADDR 855
			"00000000000000000101011010111100" , -- ADDR 856
			"00000000000000001011000011111110" , -- ADDR 857
			"00000000000000001111011000100000" , -- ADDR 858
			"00000000000000001100100000011001" , -- ADDR 859
			"00000000000000001100100100010110" , -- ADDR 860
			"00000000000000001001001100011000" , -- ADDR 861
			"00000000000000001010101010100001" , -- ADDR 862
			"00000000000000001011011111111000" , -- ADDR 863
			"00000000000000000101000001101111" , -- ADDR 864
			"00000000000000000111011000011000" , -- ADDR 865
			"00000000000000000100001011011101" , -- ADDR 866
			"00000000000000000111001110101110" , -- ADDR 867
			"00000000000000000101111101011101" , -- ADDR 868
			"00000000000000000101000101001001" , -- ADDR 869
			"00000000000000000010010011011010" , -- ADDR 870
			"00000000000000000101001000100000" , -- ADDR 871
			"00000000000000000011110011000100" , -- ADDR 872
			"00000000000000000100000100000011" , -- ADDR 873
			"00000000000000000111000001111000" , -- ADDR 874
			"00000000000000001010011111001001" , -- ADDR 875
			"00000000000000001100100110011110" , -- ADDR 876
			"00000000000000000101111001111011" , -- ADDR 877
			"00000000000000000110000000010101" , -- ADDR 878
			"00000000000000001101100111001110" , -- ADDR 879
			"00000000000000001100011100111000" , -- ADDR 880
			"00000000000000001011010100110110" , -- ADDR 881
			"00000000000000001011110101111100" , -- ADDR 882
			"00000000000000001001011001010100" , -- ADDR 883
			"00000000000000001000111000110001" , -- ADDR 884
			"00000000000000001110101011001100" , -- ADDR 885
			"00000000000000001100101111001101" , -- ADDR 886
			"00000000000000001001110111111111" , -- ADDR 887
			"00000000000000001011100010100001" , -- ADDR 888
			"00000000000000000011001011101110" , -- ADDR 889
			"00000000000000001010110011110000" , -- ADDR 890
			"00000000000000001100110001100110" , -- ADDR 891
			"00000000000000000101111000010011" , -- ADDR 892
			"00000000000000000110011111001011" , -- ADDR 893
			"00000000000000000010010000000100" , -- ADDR 894
			"00000000000000001010100010110010" , -- ADDR 895
			"00000000000000001010111010110001" , -- ADDR 896
			"00000000000000000101011000000111" , -- ADDR 897
			"00000000000000000011011011010100" , -- ADDR 898
			"00000000000000000110000100000111" , -- ADDR 899
			"00000000000000000101011101011001" , -- ADDR 900
			"00000000000000001001010010111111" , -- ADDR 901
			"00000000000000001100001111110000" , -- ADDR 902
			"00000000000000001101101001011110" , -- ADDR 903
			"00000000000000001000001101001111" , -- ADDR 904
			"00000000000000000111011110000010" , -- ADDR 905
			"00000000000000001101110100111111" , -- ADDR 906
			"00000000000000001101101111101111" , -- ADDR 907
			"00000000000000001101011101000101" , -- ADDR 908
			"00000000000000001110000011011111" , -- ADDR 909
			"00000000000000001001011000010011" , -- ADDR 910
			"00000000000000001001111100001111" , -- ADDR 911
			"00000000000000001111011000100000" , -- ADDR 912
			"00000000000000001011010000010010" , -- ADDR 913
			"00000000000000001000100011110001" , -- ADDR 914
			"00000000000000001010101110111110" , -- ADDR 915
			"00000000000000000011000001010001" , -- ADDR 916
			"00000000000000001010100000100110" , -- ADDR 917
			"00000000000000001100101111101010" , -- ADDR 918
			"00000000000000000110101010011111" , -- ADDR 919
			"00000000000000000110011010001001" , -- ADDR 920
			"00000000000000000100001101101111" , -- ADDR 921
			"00000000000000001011011000111000" , -- ADDR 922
			"00000000000000001100010001110001" , -- ADDR 923
			"00000000000000000110000111100100" , -- ADDR 924
			"00000000000000001000110011011000" , -- ADDR 925
			"00000000000000000110000111111000" , -- ADDR 926
			"00000000000000001011010010010100" , -- ADDR 927
			"00000000000000001100101100000011" , -- ADDR 928
			"00000000000000001100101111001101" , -- ADDR 929
			"00000000000000001010100010000011" , -- ADDR 930
			"00000000000000000111110100010000" , -- ADDR 931
			"00000000000000001011101110001010" , -- ADDR 932
			"00000000000000001101001111010111" , -- ADDR 933
			"00000000000000001110101111111111" , -- ADDR 934
			"00000000000000001111101000001000" , -- ADDR 935
			"00000000000000000111001111110010" , -- ADDR 936
			"00000000000000001001010011100110" , -- ADDR 937
			"00000000000000001101111000011011" , -- ADDR 938
			"00000000000000000111110100111110" , -- ADDR 939
			"00000000000000000101001011011101" , -- ADDR 940
			"00000000000000000111101001001001" , -- ADDR 941
			"00000000000000000110010111011101" , -- ADDR 942
			"00000000000000000111111100001111" , -- ADDR 943
			"00000000000000001010011000011001" , -- ADDR 944
			"00000000000000000110000110111100" , -- ADDR 945
			"00000000000000000100101000011110" , -- ADDR 946
			"00000000000000000110000010110111" , -- ADDR 947
			"00000000000000001010010011011010" , -- ADDR 948
			"00000000000000001011111101110010" , -- ADDR 949
			"00000000000000000101101000101111" , -- ADDR 950
			"00000000000000000100111100000000" , -- ADDR 951
			"00000000000000000011111010011111" , -- ADDR 952
			"00000000000000001001000000011100" , -- ADDR 953
			"00000000000000001100100011001000" , -- ADDR 954
			"00000000000000000010011101000010" , -- ADDR 955
			"00000000000000000110000000010101" , -- ADDR 956
			"00000000000000001110111001101001" , -- ADDR 957
			"00000000000000001011111010011011" , -- ADDR 958
			"00000000000000001000101000011011" , -- ADDR 959
			"00000000000000001000110010101110" , -- ADDR 960
			"00000000000000001011010010111111" , -- ADDR 961
			"00000000000000001001001011010110" , -- ADDR 962
			"00000000000000001111000111010111" , -- ADDR 963
			"00000000000000010000000011111100" , -- ADDR 964
			"00000000000000001101000111111111" , -- ADDR 965
			"00000000000000001110001111000110" , -- ADDR 966
			"00000000000000000101011101011001" , -- ADDR 967
			"00000000000000001100111101011101" , -- ADDR 968
			"00000000000000001110011101011100" , -- ADDR 969
			"00000000000000000111001011110100" , -- ADDR 970
			"00000000000000001000110011011000" , -- ADDR 971
			"00000000000000000011001101100001" , -- ADDR 972
			"00000000000000001011000001111001" , -- ADDR 973
			"00000000000000001010010111010010" , -- ADDR 974
			"00000000000000000110111000000000" , -- ADDR 975
			"00000000000000000101100111101110" , -- ADDR 976
			"00000000000000000110110101100000" , -- ADDR 977
			"00000000000000001000100010111000" , -- ADDR 978
			"00000000000000000101011001111000" , -- ADDR 979
			"00000000000000000010000000110110" , -- ADDR 980
			"00000000000000001010000100001111" , -- ADDR 981
			"00000000000000001000011010000110" , -- ADDR 982
			"00000000000000001000101000001101" , -- ADDR 983
			"00000000000000001001100011001011" , -- ADDR 984
			"00000000000000000110010111011101" , -- ADDR 985
			"00000000000000000100110110001001" , -- ADDR 986
			"00000000000000001010101110011100" , -- ADDR 987
			"00000000000000001011111011101101" , -- ADDR 988
			"00000000000000001001000000011100" , -- ADDR 989
			"00000000000000001001100010001011" , -- ADDR 990
			"00000000000000000111001111110010" , -- ADDR 991
			"00000000000000001000000011101000" , -- ADDR 992
			"00000000000000001001100010001011" , -- ADDR 993
			"00000000000000000010010000000100" , -- ADDR 994
			"00000000000000000100000101111011" , -- ADDR 995
			"00000000000000000010000110011010" , -- ADDR 996
			"00000000000000000110100100011011" , -- ADDR 997
			"00000000000000000110111001000111" , -- ADDR 998
			"00000000000000000001111101000000" , -- ADDR 999
			"00000000000000000101111010001111" , -- ADDR 1000
			"00000000000000001010011011100000" , -- ADDR 1001
			"00000000000000000001100010110101" , -- ADDR 1002
			"00000000000000000101010001010011" , -- ADDR 1003
			"00000000000000001101111011110111" , -- ADDR 1004
			"00000000000000001001011001000111" , -- ADDR 1005
			"00000000000000000100101111011000" , -- ADDR 1006
			"00000000000000000100111010000100" , -- ADDR 1007
			"00000000000000001011010011110101" , -- ADDR 1008
			"00000000000000000111110100111110" , -- ADDR 1009
			"00000000000000001101010010000110" , -- ADDR 1010
			"00000000000000010001100010111100" , -- ADDR 1011
			"00000000000000001110101000000100" , -- ADDR 1012
			"00000000000000001110111010101010" , -- ADDR 1013
			"00000000000000001001010011100110" , -- ADDR 1014
			"00000000000000001101000101100000" , -- ADDR 1015
			"00000000000000001101111100110100" , -- ADDR 1016
			"00000000000000000111010110000011" , -- ADDR 1017
			"00000000000000001001100110111101" , -- ADDR 1018
			"00000000000000000101010010000001" , -- ADDR 1019
			"00000000000000001001100110010111" , -- ADDR 1020
			"00000000000000000111111110111000" , -- ADDR 1021
			"00000000000000000111010100001111" , -- ADDR 1022
			"00000000000000000101001000001000" , -- ADDR 1023
			"00000000000000000111010000000010" , -- ADDR 1024
			"00000000000000000100111010000100" , -- ADDR 1025
			"00000000000000001001101110101010" , -- ADDR 1026
			"00000000000000000011101111000001" , -- ADDR 1027
			"00000000000000000011110010100100" , -- ADDR 1028
			"00000000000000000101010001010011" , -- ADDR 1029
			"00000000000000001000111110100010" , -- ADDR 1030
			"00000000000000000100011111010001" , -- ADDR 1031
			"00000000000000001000000011110111" , -- ADDR 1032
			"00000000000000010000100000101000" , -- ADDR 1033
			"00000000000000001101111100110100" , -- ADDR 1034
			"00000000000000001100111100101110" , -- ADDR 1035
			"00000000000000001101100001000010" , -- ADDR 1036
			"00000000000000001010100100001110" , -- ADDR 1037
			"00000000000000001010010111110101" , -- ADDR 1038
			"00000000000000000110101101111010" , -- ADDR 1039
			"00000000000000001000111101000010" , -- ADDR 1040
			"00000000000000001000001111000110" , -- ADDR 1041
			"00000000000000000101011101011001" , -- ADDR 1042
			"00000000000000000010101110101100" , -- ADDR 1043
			"00000000000000000111000111000000" , -- ADDR 1044
			"00000000000000001011011101101101" , -- ADDR 1045
			"00000000000000000110101111000010" , -- ADDR 1046
			"00000000000000000101000101001001" , -- ADDR 1047
			"00000000000000000001101000110100" , -- ADDR 1048
			"00000000000000001000110101111110" , -- ADDR 1049
			"00000000000000001010010100111001" , -- ADDR 1050
			"00000000000000000110011101101100" , -- ADDR 1051
			"00000000000000000011101110100000" , -- ADDR 1052
			"00000000000000000010111100001010" , -- ADDR 1053
			"00000000000000001101111010110001" , -- ADDR 1054
			"00000000000000001011111110000111" , -- ADDR 1055
			"00000000000000001001111100001111" , -- ADDR 1056
			"00000000000000001111110001111101" , -- ADDR 1057
			"00000000000000000111011011111111" , -- ADDR 1058
			"00000000000000000110001110010111" , -- ADDR 1059
			"00000000000000000110111111011100" , -- ADDR 1060
			"00000000000000001000001001100001" , -- ADDR 1061
			"00000000000000001010100100001110" , -- ADDR 1062
			"00000000000000000010011101000010" , -- ADDR 1063
			"00000000000000000010011111010110" , -- ADDR 1064
			"00000000000000000111100010010111" , -- ADDR 1065
			"00000000000000000101100111101110" , -- ADDR 1066
			"00000000000000001110100100100010" , -- ADDR 1067
			"00000000000000001010100100000011" , -- ADDR 1068
			"00000000000000000110010001101110" , -- ADDR 1069
			"00000000000000000110010110010000" , -- ADDR 1070
			"00000000000000001011100010100001" , -- ADDR 1071
			"00000000000000001000100001110000" , -- ADDR 1072
			"00000000000000001110001111000110" , -- ADDR 1073
			"00000000000000010001010000000101" , -- ADDR 1074
			"00000000000000001110010011100000" , -- ADDR 1075
			"00000000000000001110111011001011" , -- ADDR 1076
			"00000000000000000111111010000100" , -- ADDR 1077
			"00000000000000001101010010110100" , -- ADDR 1078
			"00000000000000001110011010011010" , -- ADDR 1079
			"00000000000000000111011011001110" , -- ADDR 1080
			"00000000000000001001011111110001" , -- ADDR 1081
			"00000000000000000100100000000111" , -- ADDR 1082
			"00000000000000001010010111010010" , -- ADDR 1083
			"00000000000000001001000101100000" , -- ADDR 1084
			"00000000000000000111010010001001" , -- ADDR 1085
			"00000000000000001001000000001110" , -- ADDR 1086
			"00000000000000000110011100110100" , -- ADDR 1087
			"00000000000000000111001011100011" , -- ADDR 1088
			"00000000000000001000010010110011" , -- ADDR 1089
			"00000000000000000110000010100011" , -- ADDR 1090
			"00000000000000000011001011101110" , -- ADDR 1091
			"00000000000000001001001001000011" , -- ADDR 1092
			"00000000000000001100101010010000" , -- ADDR 1093
			"00000000000000001001110101110111" , -- ADDR 1094
			"00000000000000001001101110000100" , -- ADDR 1095
			"00000000000000001001001011010110" , -- ADDR 1096
			"00000000000000000111110100010000" , -- ADDR 1097
			"00000000000000001000110010101110" , -- ADDR 1098
			"00000000000000000010010000000100" , -- ADDR 1099
			"00000000000000000100101010100001" , -- ADDR 1100
			"00000000000000000011110111000011" , -- ADDR 1101
			"00000000000000000101000001101111" , -- ADDR 1102
			"00000000000000000100111010011101" , -- ADDR 1103
			"00000000000000000010011100010000" , -- ADDR 1104
			"00000000000000000110101101000011" , -- ADDR 1105
			"00000000000000001101100001000010" , -- ADDR 1106
			"00000000000000001110111111011000" , -- ADDR 1107
			"00000000000000000100100000000111" , -- ADDR 1108
			"00000000000000000110000110111100" , -- ADDR 1109
			"00000000000000000011011001101000" , -- ADDR 1110
			"00000000000000001010000011101011" , -- ADDR 1111
			"00000000000000001000111101000010" , -- ADDR 1112
			"00000000000000000110000110101000" , -- ADDR 1113
			"00000000000000010000100011011001" , -- ADDR 1114
			"00000000000000000100000101111011" , -- ADDR 1115
			"00000000000000000001101101011000" , -- ADDR 1116
			"00000000000000000111110111001010" , -- ADDR 1117
			"00000000000000000111011011001110" , -- ADDR 1118
			"00000000000000001100000111111011" , -- ADDR 1119
			"00000000000000000100011010111111" , -- ADDR 1120
			"00000000000000000111000001111000" , -- ADDR 1121
			"00000000000000001000010011010000" , -- ADDR 1122
			"00000000000000000111010101000001" , -- ADDR 1123
			"00000000000000001000110011011000" , -- ADDR 1124
			"00000000000000000111100100101000" , -- ADDR 1125
			"00000000000000000011111011111101" , -- ADDR 1126
			"00000000000000000100011010111111" , -- ADDR 1127
			"00000000000000001111001011011001" , -- ADDR 1128
			"00000000000000001101000011001011" , -- ADDR 1129
			"00000000000000001011010000111101" , -- ADDR 1130
			"00000000000000001111101000001000" , -- ADDR 1131
			"00000000000000001000110000000111" , -- ADDR 1132
			"00000000000000000111110001010100" , -- ADDR 1133
			"00000000000000000111001110101110" , -- ADDR 1134
			"00000000000000001000110010101110" , -- ADDR 1135
			"00000000000000001010010011001110" , -- ADDR 1136
			"00000000000000000011011001101000" , -- ADDR 1137
			"00000000000000000001100100000011" , -- ADDR 1138
			"00000000000000000111110000100100" , -- ADDR 1139
			"00000000000000000001011111000011" , -- ADDR 1140
			"00000000000000001100011001110100" , -- ADDR 1141
			"00000000000000000111111111110101" , -- ADDR 1142
			"00000000000000001011101111011110" , -- ADDR 1143
			"00000000000000010011101011100010" , -- ADDR 1144
			"00000000000000010000111100110010" , -- ADDR 1145
			"00000000000000010000010110111111" , -- ADDR 1146
			"00000000000000001101111010110001" , -- ADDR 1147
			"00000000000000001110000101011001" , -- ADDR 1148
			"00000000000000001110000110101111" , -- ADDR 1149
			"00000000000000001001011000010011" , -- ADDR 1150
			"00000000000000001011110010001110" , -- ADDR 1151
			"00000000000000001001001111011111" , -- ADDR 1152
			"00000000000000001001001101000000" , -- ADDR 1153
			"00000000000000000110100000111011" , -- ADDR 1154
			"00000000000000001001100111110000" , -- ADDR 1155
			"00000000000000001101101111101111" , -- ADDR 1156
			"00000000000000001001011001000111" , -- ADDR 1157
			"00000000000000001101001110000100" , -- ADDR 1158
			"00000000000000010100111010000001" , -- ADDR 1159
			"00000000000000010010001000001010" , -- ADDR 1160
			"00000000000000010001101011100110" , -- ADDR 1161
			"00000000000000001110001101100111" , -- ADDR 1162
			"00000000000000001111011100110101" , -- ADDR 1163
			"00000000000000001111100011001111" , -- ADDR 1164
			"00000000000000001010100010000011" , -- ADDR 1165
			"00000000000000001100111100101110" , -- ADDR 1166
			"00000000000000001001111000110001" , -- ADDR 1167
			"00000000000000001010101010001010" , -- ADDR 1168
			"00000000000000000111111111110101" , -- ADDR 1169
			"00000000000000001010101110011100" , -- ADDR 1170
			"00000000000000000100011111010001" , -- ADDR 1171
			"00000000000000000110110011110101" , -- ADDR 1172
			"00000000000000000111101010011001" , -- ADDR 1173
			"00000000000000000101100000100001" , -- ADDR 1174
			"00000000000000000011111110010111" , -- ADDR 1175
			"00000000000000001100001100001010" , -- ADDR 1176
			"00000000000000000001110001110000" , -- ADDR 1177
			"00000000000000000011011001000100" , -- ADDR 1178
			"00000000000000000100001001101000" , -- ADDR 1179
			"00000000000000000010111110101111" , -- ADDR 1180
			"00000000000000001000001111000110" , -- ADDR 1181
			"00000000000000000100001011000000" , -- ADDR 1182
			"00000000000000000110111010001110" , -- ADDR 1183
			"00000000000000000100011010111111" , -- ADDR 1184
			"00000000000000000101111101011101" , -- ADDR 1185
			"00000000000000001100000011111110" , -- ADDR 1186
			"00000000000000001001100110111101" , -- ADDR 1187
			"00000000000000001000011101011111" , -- ADDR 1188
			"00000000000000001100000011111110" , -- ADDR 1189
			"00000000000000000110000110101000" , -- ADDR 1190
			"00000000000000000110010001101110" , -- ADDR 1191
			"00000000000000000011010100100001" , -- ADDR 1192
			"00000000000000000100111100000000" , -- ADDR 1193
			"00000000000000000110111001111100" , -- ADDR 1194
			"00000000000000000001110111000000" , -- ADDR 1195
			"00000000000000000010101110101100" , -- ADDR 1196
			"00000000000000000011110111000011" , -- ADDR 1197
			"00000000000000001101010111011001" , -- ADDR 1198
			"00000000000000001011111110010001" , -- ADDR 1199
			"00000000000000001001010110111000" , -- ADDR 1200
			"00000000000000010001110011010110" , -- ADDR 1201
			"00000000000000000111000101001000" , -- ADDR 1202
			"00000000000000000101000010001000" , -- ADDR 1203
			"00000000000000001000110100011101" , -- ADDR 1204
			"00000000000000001001010001111101" , -- ADDR 1205
			"00000000000000001100110100010010" , -- ADDR 1206
			"00000000000000000100001010000101" , -- ADDR 1207
			"00000000000000000101011010111100" , -- ADDR 1208
			"00000000000000001001010110010000" , -- ADDR 1209
			"00000000000000000010111100110011" , -- ADDR 1210
			"00000000000000000100000001101100" , -- ADDR 1211
			"00000000000000001110001010010000" , -- ADDR 1212
			"00000000000000000110011111001011" , -- ADDR 1213
			"00000000000000001000010110111010" , -- ADDR 1214
			"00000000000000001010011010001110" , -- ADDR 1215
			"00000000000000001000000000100010" , -- ADDR 1216
			"00000000000000001100111010111100" , -- ADDR 1217
			"00000000000000001011110010101101" , -- ADDR 1218
			"00000000000000001110100100100010" , -- ADDR 1219
			"00000000000000001010010011011010" , -- ADDR 1220
			"00000000000000000011001011101110" , -- ADDR 1221
			"00000000000000001011100010100001" , -- ADDR 1222
			"00000000000000000100111010000100" , -- ADDR 1223
			"00000000000000000111010010001001" , -- ADDR 1224
			"00000000000000000111100110001001" , -- ADDR 1225
			"00000000000000000101001011011101" , -- ADDR 1226
			"00000000000000001001111110010101" , -- ADDR 1227
			"00000000000000001001101010001000" , -- ADDR 1228
			"00000000000000001100001111110000" , -- ADDR 1229
			"00000000000000000111011100010000" , -- ADDR 1230
			"00000000000000001101110000000001" , -- ADDR 1231
			"00000000000000000010100000111000" , -- ADDR 1232
			"00000000000000000100011001010000" , -- ADDR 1233
			"00000000000000000111100100101000" , -- ADDR 1234
			"00000000000000000101011101011001" , -- ADDR 1235
			"00000000000000001011000001111001" , -- ADDR 1236
			"00000000000000000111111011000010" , -- ADDR 1237
			"00000000000000001010110010101100" , -- ADDR 1238
			"00000000000000000111101001011001" , -- ADDR 1239
			"00000000000000001101011011100001" , -- ADDR 1240
			"00000000000000001111100101000100" , -- ADDR 1241
			"00000000000000001000111110111101" , -- ADDR 1242
			"00000000000000001001001101101000" , -- ADDR 1243
			"00000000000000000101010110101100" , -- ADDR 1244
			"00000000000000001101101100010000" , -- ADDR 1245
			"00000000000000001110000101101010" , -- ADDR 1246
			"00000000000000001000011101011111" , -- ADDR 1247
			"00000000000000000010100000111000" , -- ADDR 1248
			"00000000000000000101111000010011" , -- ADDR 1249
			"00000000000000000100010100111000" , -- ADDR 1250
			"00000000000000001001110101110111" , -- ADDR 1251
			"00000000000000000101011010111100" , -- ADDR 1252
			"00000000000000001000010100001011" , -- ADDR 1253
			"00000000000000000110000110101000" , -- ADDR 1254
			"00000000000000000111010010001001" , -- ADDR 1255
			"00000000000000000110010111011101" , -- ADDR 1256
			"00000000000000001011100000010111" , -- ADDR 1257
			"00000000000000000100111010011101" , -- ADDR 1258
			"00000000000000000111110010100010" , -- ADDR 1259
			"00000000000000000111101001011001" , -- ADDR 1260
			"00000000000000000010011010101011" , -- ADDR 1261
			"00000000000000000100010000111000" , -- ADDR 1262
			"00000000000000000100101111011000" , -- ADDR 1263
			"00000000000000000101111000010011" , -- ADDR 1264
			"00000000000000000000100010111100" , -- ADDR 1265
			"00000000000000000101100111011000" , -- ADDR 1266
			"00000000000000000101101100110001" , -- ADDR 1267
			"00000000000000000111101010101001" , -- ADDR 1268
			"00000000000000000010010011011010" , -- ADDR 1269
			"00000000000000001000101010001100" , -- ADDR 1270
			"00000000000000001000110000000111" , -- ADDR 1271
			"00000000000000000011110111000011" , -- ADDR 1272
			"00000000000000000010111100001010" , -- ADDR 1273
			"00000000000000000101010010000001" , -- ADDR 1274
			"00000000000000000110011000111101" , -- ADDR 1275
			"00000000000000000000000000000000" , -- ADDR 1276
			"00000000000000000000000000000000" , -- ADDR 1277
			"00000000000000000000000000000000" , -- ADDR 1278
			"00000000000000000000000000000000" , -- ADDR 1279
			"00000000000000000000000000000000" , -- ADDR 1280
			"00000000000000000000000000000000" , -- ADDR 1281
			"00000000000000000000000000000000" , -- ADDR 1282
			"00000000000000000000000000000000" , -- ADDR 1283
			"00000000000000000000000000000000" , -- ADDR 1284
			"00000000000000000000000000000000" , -- ADDR 1285
			"00000000000000000000000000000000" , -- ADDR 1286
			"00000000000000000000000000000000" , -- ADDR 1287
			"00000000000000000000000000000000" , -- ADDR 1288
			"00000000000000000000000000000000" , -- ADDR 1289
			"00000000000000000000000000000000" , -- ADDR 1290
			"00000000000000000000000000000000" , -- ADDR 1291
			"00000000000000000000000000000000" , -- ADDR 1292
			"00000000000000000000000000000000" , -- ADDR 1293
			"00000000000000000000000000000000" , -- ADDR 1294
			"00000000000000000000000000000000" , -- ADDR 1295
			"00000000000000000000000000000000" , -- ADDR 1296
			"00000000000000000000000000000000" , -- ADDR 1297
			"00000000000000000000000000000000" , -- ADDR 1298
			"00000000000000000000000000000000" , -- ADDR 1299
			"00000000000000000000000000000000" , -- ADDR 1300
			"00000000000000000000000000000000" , -- ADDR 1301
			"00000000000000000000000000000000" , -- ADDR 1302
			"00000000000000000000000000000000" , -- ADDR 1303
			"00000000000000000000000000000000" , -- ADDR 1304
			"00000000000000000000000000000000" , -- ADDR 1305
			"00000000000000000000000000000000" , -- ADDR 1306
			"00000000000000000000000000000000" , -- ADDR 1307
			"00000000000000000000000000000000" , -- ADDR 1308
			"00000000000000000000000000000000" , -- ADDR 1309
			"00000000000000000000000000000000" , -- ADDR 1310
			"00000000000000000000000000000000" , -- ADDR 1311
			"00000000000000000000000000000000" , -- ADDR 1312
			"00000000000000000000000000000000" , -- ADDR 1313
			"00000000000000000000000000000000" , -- ADDR 1314
			"00000000000000000000000000000000" , -- ADDR 1315
			"00000000000000000000000000000000" , -- ADDR 1316
			"00000000000000000000000000000000" , -- ADDR 1317
			"00000000000000000000000000000000" , -- ADDR 1318
			"00000000000000000000000000000000" , -- ADDR 1319
			"00000000000000000000000000000000" , -- ADDR 1320
			"00000000000000000000000000000000" , -- ADDR 1321
			"00000000000000000000000000000000" , -- ADDR 1322
			"00000000000000000000000000000000" , -- ADDR 1323
			"00000000000000000000000000000000" , -- ADDR 1324
			"00000000000000000000000000000000" , -- ADDR 1325
			"00000000000000000000000000000000" , -- ADDR 1326
			"00000000000000000000000000000000" , -- ADDR 1327
			"00000000000000000000000000000000" , -- ADDR 1328
			"00000000000000000000000000000000" , -- ADDR 1329
			"00000000000000000000000000000000" , -- ADDR 1330
			"00000000000000000000000000000000" , -- ADDR 1331
			"00000000000000000000000000000000" , -- ADDR 1332
			"00000000000000000000000000000000" , -- ADDR 1333
			"00000000000000000000000000000000" , -- ADDR 1334
			"00000000000000000000000000000000" , -- ADDR 1335
			"00000000000000000000000000000000" , -- ADDR 1336
			"00000000000000000000000000000000" , -- ADDR 1337
			"00000000000000000000000000000000" , -- ADDR 1338
			"00000000000000000000000000000000" , -- ADDR 1339
			"00000000000000000000000000000000" , -- ADDR 1340
			"00000000000000000000000000000000" , -- ADDR 1341
			"00000000000000000000000000000000" , -- ADDR 1342
			"00000000000000000000000000000000" , -- ADDR 1343
			"00000000000000000000000000000000" , -- ADDR 1344
			"00000000000000000000000000000000" , -- ADDR 1345
			"00000000000000000000000000000000" , -- ADDR 1346
			"00000000000000000000000000000000" , -- ADDR 1347
			"00000000000000000000000000000000" , -- ADDR 1348
			"00000000000000000000000000000000" , -- ADDR 1349
			"00000000000000000000000000000000" , -- ADDR 1350
			"00000000000000000000000000000000" , -- ADDR 1351
			"00000000000000000000000000000000" , -- ADDR 1352
			"00000000000000000000000000000000" , -- ADDR 1353
			"00000000000000000000000000000000" , -- ADDR 1354
			"00000000000000000000000000000000" , -- ADDR 1355
			"00000000000000000000000000000000" , -- ADDR 1356
			"00000000000000000000000000000000" , -- ADDR 1357
			"00000000000000000000000000000000" , -- ADDR 1358
			"00000000000000000000000000000000" , -- ADDR 1359
			"00000000000000000000000000000000" , -- ADDR 1360
			"00000000000000000000000000000000" , -- ADDR 1361
			"00000000000000000000000000000000" , -- ADDR 1362
			"00000000000000000000000000000000" , -- ADDR 1363
			"00000000000000000000000000000000" , -- ADDR 1364
			"00000000000000000000000000000000" , -- ADDR 1365
			"00000000000000000000000000000000" , -- ADDR 1366
			"00000000000000000000000000000000" , -- ADDR 1367
			"00000000000000000000000000000000" , -- ADDR 1368
			"00000000000000000000000000000000" , -- ADDR 1369
			"00000000000000000000000000000000" , -- ADDR 1370
			"00000000000000000000000000000000" , -- ADDR 1371
			"00000000000000000000000000000000" , -- ADDR 1372
			"00000000000000000000000000000000" , -- ADDR 1373
			"00000000000000000000000000000000" , -- ADDR 1374
			"00000000000000000000000000000000" , -- ADDR 1375
			"00000000000000000000000000000000" , -- ADDR 1376
			"00000000000000000000000000000000" , -- ADDR 1377
			"00000000000000000000000000000000" , -- ADDR 1378
			"00000000000000000000000000000000" , -- ADDR 1379
			"00000000000000000000000000000000" , -- ADDR 1380
			"00000000000000000000000000000000" , -- ADDR 1381
			"00000000000000000000000000000000" , -- ADDR 1382
			"00000000000000000000000000000000" , -- ADDR 1383
			"00000000000000000000000000000000" , -- ADDR 1384
			"00000000000000000000000000000000" , -- ADDR 1385
			"00000000000000000000000000000000" , -- ADDR 1386
			"00000000000000000000000000000000" , -- ADDR 1387
			"00000000000000000000000000000000" , -- ADDR 1388
			"00000000000000000000000000000000" , -- ADDR 1389
			"00000000000000000000000000000000" , -- ADDR 1390
			"00000000000000000000000000000000" , -- ADDR 1391
			"00000000000000000000000000000000" , -- ADDR 1392
			"00000000000000000000000000000000" , -- ADDR 1393
			"00000000000000000000000000000000" , -- ADDR 1394
			"00000000000000000000000000000000" , -- ADDR 1395
			"00000000000000000000000000000000" , -- ADDR 1396
			"00000000000000000000000000000000" , -- ADDR 1397
			"00000000000000000000000000000000" , -- ADDR 1398
			"00000000000000000000000000000000" , -- ADDR 1399
			"00000000000000000000000000000000" , -- ADDR 1400
			"00000000000000000000000000000000" , -- ADDR 1401
			"00000000000000000000000000000000" , -- ADDR 1402
			"00000000000000000000000000000000" , -- ADDR 1403
			"00000000000000000000000000000000" , -- ADDR 1404
			"00000000000000000000000000000000" , -- ADDR 1405
			"00000000000000000000000000000000" , -- ADDR 1406
			"00000000000000000000000000000000" , -- ADDR 1407
			"00000000000000000000000000000000" , -- ADDR 1408
			"00000000000000000000000000000000" , -- ADDR 1409
			"00000000000000000000000000000000" , -- ADDR 1410
			"00000000000000000000000000000000" , -- ADDR 1411
			"00000000000000000000000000000000" , -- ADDR 1412
			"00000000000000000000000000000000" , -- ADDR 1413
			"00000000000000000000000000000000" , -- ADDR 1414
			"00000000000000000000000000000000" , -- ADDR 1415
			"00000000000000000000000000000000" , -- ADDR 1416
			"00000000000000000000000000000000" , -- ADDR 1417
			"00000000000000000000000000000000" , -- ADDR 1418
			"00000000000000000000000000000000" , -- ADDR 1419
			"00000000000000000000000000000000" , -- ADDR 1420
			"00000000000000000000000000000000" , -- ADDR 1421
			"00000000000000000000000000000000" , -- ADDR 1422
			"00000000000000000000000000000000" , -- ADDR 1423
			"00000000000000000000000000000000" , -- ADDR 1424
			"00000000000000000000000000000000" , -- ADDR 1425
			"00000000000000000000000000000000" , -- ADDR 1426
			"00000000000000000000000000000000" , -- ADDR 1427
			"00000000000000000000000000000000" , -- ADDR 1428
			"00000000000000000000000000000000" , -- ADDR 1429
			"00000000000000000000000000000000" , -- ADDR 1430
			"00000000000000000000000000000000" , -- ADDR 1431
			"00000000000000000000000000000000" , -- ADDR 1432
			"00000000000000000000000000000000" , -- ADDR 1433
			"00000000000000000000000000000000" , -- ADDR 1434
			"00000000000000000000000000000000" , -- ADDR 1435
			"00000000000000000000000000000000" , -- ADDR 1436
			"00000000000000000000000000000000" , -- ADDR 1437
			"00000000000000000000000000000000" , -- ADDR 1438
			"00000000000000000000000000000000" , -- ADDR 1439
			"00000000000000000000000000000000" , -- ADDR 1440
			"00000000000000000000000000000000" , -- ADDR 1441
			"00000000000000000000000000000000" , -- ADDR 1442
			"00000000000000000000000000000000" , -- ADDR 1443
			"00000000000000000000000000000000" , -- ADDR 1444
			"00000000000000000000000000000000" , -- ADDR 1445
			"00000000000000000000000000000000" , -- ADDR 1446
			"00000000000000000000000000000000" , -- ADDR 1447
			"00000000000000000000000000000000" , -- ADDR 1448
			"00000000000000000000000000000000" , -- ADDR 1449
			"00000000000000000000000000000000" , -- ADDR 1450
			"00000000000000000000000000000000" , -- ADDR 1451
			"00000000000000000000000000000000" , -- ADDR 1452
			"00000000000000000000000000000000" , -- ADDR 1453
			"00000000000000000000000000000000" , -- ADDR 1454
			"00000000000000000000000000000000" , -- ADDR 1455
			"00000000000000000000000000000000" , -- ADDR 1456
			"00000000000000000000000000000000" , -- ADDR 1457
			"00000000000000000000000000000000" , -- ADDR 1458
			"00000000000000000000000000000000" , -- ADDR 1459
			"00000000000000000000000000000000" , -- ADDR 1460
			"00000000000000000000000000000000" , -- ADDR 1461
			"00000000000000000000000000000000" , -- ADDR 1462
			"00000000000000000000000000000000" , -- ADDR 1463
			"00000000000000000000000000000000" , -- ADDR 1464
			"00000000000000000000000000000000" , -- ADDR 1465
			"00000000000000000000000000000000" , -- ADDR 1466
			"00000000000000000000000000000000" , -- ADDR 1467
			"00000000000000000000000000000000" , -- ADDR 1468
			"00000000000000000000000000000000" , -- ADDR 1469
			"00000000000000000000000000000000" , -- ADDR 1470
			"00000000000000000000000000000000" , -- ADDR 1471
			"00000000000000000000000000000000" , -- ADDR 1472
			"00000000000000000000000000000000" , -- ADDR 1473
			"00000000000000000000000000000000" , -- ADDR 1474
			"00000000000000000000000000000000" , -- ADDR 1475
			"00000000000000000000000000000000" , -- ADDR 1476
			"00000000000000000000000000000000" , -- ADDR 1477
			"00000000000000000000000000000000" , -- ADDR 1478
			"00000000000000000000000000000000" , -- ADDR 1479
			"00000000000000000000000000000000" , -- ADDR 1480
			"00000000000000000000000000000000" , -- ADDR 1481
			"00000000000000000000000000000000" , -- ADDR 1482
			"00000000000000000000000000000000" , -- ADDR 1483
			"00000000000000000000000000000000" , -- ADDR 1484
			"00000000000000000000000000000000" , -- ADDR 1485
			"00000000000000000000000000000000" , -- ADDR 1486
			"00000000000000000000000000000000" , -- ADDR 1487
			"00000000000000000000000000000000" , -- ADDR 1488
			"00000000000000000000000000000000" , -- ADDR 1489
			"00000000000000000000000000000000" , -- ADDR 1490
			"00000000000000000000000000000000" , -- ADDR 1491
			"00000000000000000000000000000000" , -- ADDR 1492
			"00000000000000000000000000000000" , -- ADDR 1493
			"00000000000000000000000000000000" , -- ADDR 1494
			"00000000000000000000000000000000" , -- ADDR 1495
			"00000000000000000000000000000000" , -- ADDR 1496
			"00000000000000000000000000000000" , -- ADDR 1497
			"00000000000000000000000000000000" , -- ADDR 1498
			"00000000000000000000000000000000" , -- ADDR 1499
			"00000000000000000000000000000000" , -- ADDR 1500
			"00000000000000000000000000000000" , -- ADDR 1501
			"00000000000000000000000000000000" , -- ADDR 1502
			"00000000000000000000000000000000" , -- ADDR 1503
			"00000000000000000000000000000000" , -- ADDR 1504
			"00000000000000000000000000000000" , -- ADDR 1505
			"00000000000000000000000000000000" , -- ADDR 1506
			"00000000000000000000000000000000" , -- ADDR 1507
			"00000000000000000000000000000000" , -- ADDR 1508
			"00000000000000000000000000000000" , -- ADDR 1509
			"00000000000000000000000000000000" , -- ADDR 1510
			"00000000000000000000000000000000" , -- ADDR 1511
			"00000000000000000000000000000000" , -- ADDR 1512
			"00000000000000000000000000000000" , -- ADDR 1513
			"00000000000000000000000000000000" , -- ADDR 1514
			"00000000000000000000000000000000" , -- ADDR 1515
			"00000000000000000000000000000000" , -- ADDR 1516
			"00000000000000000000000000000000" , -- ADDR 1517
			"00000000000000000000000000000000" , -- ADDR 1518
			"00000000000000000000000000000000" , -- ADDR 1519
			"00000000000000000000000000000000" , -- ADDR 1520
			"00000000000000000000000000000000" , -- ADDR 1521
			"00000000000000000000000000000000" , -- ADDR 1522
			"00000000000000000000000000000000" , -- ADDR 1523
			"00000000000000000000000000000000" , -- ADDR 1524
			"00000000000000000000000000000000" , -- ADDR 1525
			"00000000000000000000000000000000" , -- ADDR 1526
			"00000000000000000000000000000000" , -- ADDR 1527
			"00000000000000000000000000000000" , -- ADDR 1528
			"00000000000000000000000000000000" , -- ADDR 1529
			"00000000000000000000000000000000" , -- ADDR 1530
			"00000000000000000000000000000000" , -- ADDR 1531
			"00000000000000000000000000000000" , -- ADDR 1532
			"00000000000000000000000000000000" , -- ADDR 1533
			"00000000000000000000000000000000" , -- ADDR 1534
			"00000000000000000000000000000000" , -- ADDR 1535
			"00000000000000000000000000000000" , -- ADDR 1536
			"00000000000000000000000000000000" , -- ADDR 1537
			"00000000000000000000000000000000" , -- ADDR 1538
			"00000000000000000000000000000000" , -- ADDR 1539
			"00000000000000000000000000000000" , -- ADDR 1540
			"00000000000000000000000000000000" , -- ADDR 1541
			"00000000000000000000000000000000" , -- ADDR 1542
			"00000000000000000000000000000000" , -- ADDR 1543
			"00000000000000000000000000000000" , -- ADDR 1544
			"00000000000000000000000000000000" , -- ADDR 1545
			"00000000000000000000000000000000" , -- ADDR 1546
			"00000000000000000000000000000000" , -- ADDR 1547
			"00000000000000000000000000000000" , -- ADDR 1548
			"00000000000000000000000000000000" , -- ADDR 1549
			"00000000000000000000000000000000" , -- ADDR 1550
			"00000000000000000000000000000000" , -- ADDR 1551
			"00000000000000000000000000000000" , -- ADDR 1552
			"00000000000000000000000000000000" , -- ADDR 1553
			"00000000000000000000000000000000" , -- ADDR 1554
			"00000000000000000000000000000000" , -- ADDR 1555
			"00000000000000000000000000000000" , -- ADDR 1556
			"00000000000000000000000000000000" , -- ADDR 1557
			"00000000000000000000000000000000" , -- ADDR 1558
			"00000000000000000000000000000000" , -- ADDR 1559
			"00000000000000000000000000000000" , -- ADDR 1560
			"00000000000000000000000000000000" , -- ADDR 1561
			"00000000000000000000000000000000" , -- ADDR 1562
			"00000000000000000000000000000000" , -- ADDR 1563
			"00000000000000000000000000000000" , -- ADDR 1564
			"00000000000000000000000000000000" , -- ADDR 1565
			"00000000000000000000000000000000" , -- ADDR 1566
			"00000000000000000000000000000000" , -- ADDR 1567
			"00000000000000000000000000000000" , -- ADDR 1568
			"00000000000000000000000000000000" , -- ADDR 1569
			"00000000000000000000000000000000" , -- ADDR 1570
			"00000000000000000000000000000000" , -- ADDR 1571
			"00000000000000000000000000000000" , -- ADDR 1572
			"00000000000000000000000000000000" , -- ADDR 1573
			"00000000000000000000000000000000" , -- ADDR 1574
			"00000000000000000000000000000000" , -- ADDR 1575
			"00000000000000000000000000000000" , -- ADDR 1576
			"00000000000000000000000000000000" , -- ADDR 1577
			"00000000000000000000000000000000" , -- ADDR 1578
			"00000000000000000000000000000000" , -- ADDR 1579
			"00000000000000000000000000000000" , -- ADDR 1580
			"00000000000000000000000000000000" , -- ADDR 1581
			"00000000000000000000000000000000" , -- ADDR 1582
			"00000000000000000000000000000000" , -- ADDR 1583
			"00000000000000000000000000000000" , -- ADDR 1584
			"00000000000000000000000000000000" , -- ADDR 1585
			"00000000000000000000000000000000" , -- ADDR 1586
			"00000000000000000000000000000000" , -- ADDR 1587
			"00000000000000000000000000000000" , -- ADDR 1588
			"00000000000000000000000000000000" , -- ADDR 1589
			"00000000000000000000000000000000" , -- ADDR 1590
			"00000000000000000000000000000000" , -- ADDR 1591
			"00000000000000000000000000000000" , -- ADDR 1592
			"00000000000000000000000000000000" , -- ADDR 1593
			"00000000000000000000000000000000" , -- ADDR 1594
			"00000000000000000000000000000000" , -- ADDR 1595
			"00000000000000000000000000000000" , -- ADDR 1596
			"00000000000000000000000000000000" , -- ADDR 1597
			"00000000000000000000000000000000" , -- ADDR 1598
			"00000000000000000000000000000000" , -- ADDR 1599
			"00000000000000000000000000000000" , -- ADDR 1600
			"00000000000000000000000000000000" , -- ADDR 1601
			"00000000000000000000000000000000" , -- ADDR 1602
			"00000000000000000000000000000000" , -- ADDR 1603
			"00000000000000000000000000000000" , -- ADDR 1604
			"00000000000000000000000000000000" , -- ADDR 1605
			"00000000000000000000000000000000" , -- ADDR 1606
			"00000000000000000000000000000000" , -- ADDR 1607
			"00000000000000000000000000000000" , -- ADDR 1608
			"00000000000000000000000000000000" , -- ADDR 1609
			"00000000000000000000000000000000" , -- ADDR 1610
			"00000000000000000000000000000000" , -- ADDR 1611
			"00000000000000000000000000000000" , -- ADDR 1612
			"00000000000000000000000000000000" , -- ADDR 1613
			"00000000000000000000000000000000" , -- ADDR 1614
			"00000000000000000000000000000000" , -- ADDR 1615
			"00000000000000000000000000000000" , -- ADDR 1616
			"00000000000000000000000000000000" , -- ADDR 1617
			"00000000000000000000000000000000" , -- ADDR 1618
			"00000000000000000000000000000000" , -- ADDR 1619
			"00000000000000000000000000000000" , -- ADDR 1620
			"00000000000000000000000000000000" , -- ADDR 1621
			"00000000000000000000000000000000" , -- ADDR 1622
			"00000000000000000000000000000000" , -- ADDR 1623
			"00000000000000000000000000000000" , -- ADDR 1624
			"00000000000000000000000000000000" , -- ADDR 1625
			"00000000000000000000000000000000" , -- ADDR 1626
			"00000000000000000000000000000000" , -- ADDR 1627
			"00000000000000000000000000000000" , -- ADDR 1628
			"00000000000000000000000000000000" , -- ADDR 1629
			"00000000000000000000000000000000" , -- ADDR 1630
			"00000000000000000000000000000000" , -- ADDR 1631
			"00000000000000000000000000000000" , -- ADDR 1632
			"00000000000000000000000000000000" , -- ADDR 1633
			"00000000000000000000000000000000" , -- ADDR 1634
			"00000000000000000000000000000000" , -- ADDR 1635
			"00000000000000000000000000000000" , -- ADDR 1636
			"00000000000000000000000000000000" , -- ADDR 1637
			"00000000000000000000000000000000" , -- ADDR 1638
			"00000000000000000000000000000000" , -- ADDR 1639
			"00000000000000000000000000000000" , -- ADDR 1640
			"00000000000000000000000000000000" , -- ADDR 1641
			"00000000000000000000000000000000" , -- ADDR 1642
			"00000000000000000000000000000000" , -- ADDR 1643
			"00000000000000000000000000000000" , -- ADDR 1644
			"00000000000000000000000000000000" , -- ADDR 1645
			"00000000000000000000000000000000" , -- ADDR 1646
			"00000000000000000000000000000000" , -- ADDR 1647
			"00000000000000000000000000000000" , -- ADDR 1648
			"00000000000000000000000000000000" , -- ADDR 1649
			"00000000000000000000000000000000" , -- ADDR 1650
			"00000000000000000000000000000000" , -- ADDR 1651
			"00000000000000000000000000000000" , -- ADDR 1652
			"00000000000000000000000000000000" , -- ADDR 1653
			"00000000000000000000000000000000" , -- ADDR 1654
			"00000000000000000000000000000000" , -- ADDR 1655
			"00000000000000000000000000000000" , -- ADDR 1656
			"00000000000000000000000000000000" , -- ADDR 1657
			"00000000000000000000000000000000" , -- ADDR 1658
			"00000000000000000000000000000000" , -- ADDR 1659
			"00000000000000000000000000000000" , -- ADDR 1660
			"00000000000000000000000000000000" , -- ADDR 1661
			"00000000000000000000000000000000" , -- ADDR 1662
			"00000000000000000000000000000000" , -- ADDR 1663
			"00000000000000000000000000000000" , -- ADDR 1664
			"00000000000000000000000000000000" , -- ADDR 1665
			"00000000000000000000000000000000" , -- ADDR 1666
			"00000000000000000000000000000000" , -- ADDR 1667
			"00000000000000000000000000000000" , -- ADDR 1668
			"00000000000000000000000000000000" , -- ADDR 1669
			"00000000000000000000000000000000" , -- ADDR 1670
			"00000000000000000000000000000000" , -- ADDR 1671
			"00000000000000000000000000000000" , -- ADDR 1672
			"00000000000000000000000000000000" , -- ADDR 1673
			"00000000000000000000000000000000" , -- ADDR 1674
			"00000000000000000000000000000000" , -- ADDR 1675
			"00000000000000000000000000000000" , -- ADDR 1676
			"00000000000000000000000000000000" , -- ADDR 1677
			"00000000000000000000000000000000" , -- ADDR 1678
			"00000000000000000000000000000000" , -- ADDR 1679
			"00000000000000000000000000000000" , -- ADDR 1680
			"00000000000000000000000000000000" , -- ADDR 1681
			"00000000000000000000000000000000" , -- ADDR 1682
			"00000000000000000000000000000000" , -- ADDR 1683
			"00000000000000000000000000000000" , -- ADDR 1684
			"00000000000000000000000000000000" , -- ADDR 1685
			"00000000000000000000000000000000" , -- ADDR 1686
			"00000000000000000000000000000000" , -- ADDR 1687
			"00000000000000000000000000000000" , -- ADDR 1688
			"00000000000000000000000000000000" , -- ADDR 1689
			"00000000000000000000000000000000" , -- ADDR 1690
			"00000000000000000000000000000000" , -- ADDR 1691
			"00000000000000000000000000000000" , -- ADDR 1692
			"00000000000000000000000000000000" , -- ADDR 1693
			"00000000000000000000000000000000" , -- ADDR 1694
			"00000000000000000000000000000000" , -- ADDR 1695
			"00000000000000000000000000000000" , -- ADDR 1696
			"00000000000000000000000000000000" , -- ADDR 1697
			"00000000000000000000000000000000" , -- ADDR 1698
			"00000000000000000000000000000000" , -- ADDR 1699
			"00000000000000000000000000000000" , -- ADDR 1700
			"00000000000000000000000000000000" , -- ADDR 1701
			"00000000000000000000000000000000" , -- ADDR 1702
			"00000000000000000000000000000000" , -- ADDR 1703
			"00000000000000000000000000000000" , -- ADDR 1704
			"00000000000000000000000000000000" , -- ADDR 1705
			"00000000000000000000000000000000" , -- ADDR 1706
			"00000000000000000000000000000000" , -- ADDR 1707
			"00000000000000000000000000000000" , -- ADDR 1708
			"00000000000000000000000000000000" , -- ADDR 1709
			"00000000000000000000000000000000" , -- ADDR 1710
			"00000000000000000000000000000000" , -- ADDR 1711
			"00000000000000000000000000000000" , -- ADDR 1712
			"00000000000000000000000000000000" , -- ADDR 1713
			"00000000000000000000000000000000" , -- ADDR 1714
			"00000000000000000000000000000000" , -- ADDR 1715
			"00000000000000000000000000000000" , -- ADDR 1716
			"00000000000000000000000000000000" , -- ADDR 1717
			"00000000000000000000000000000000" , -- ADDR 1718
			"00000000000000000000000000000000" , -- ADDR 1719
			"00000000000000000000000000000000" , -- ADDR 1720
			"00000000000000000000000000000000" , -- ADDR 1721
			"00000000000000000000000000000000" , -- ADDR 1722
			"00000000000000000000000000000000" , -- ADDR 1723
			"00000000000000000000000000000000" , -- ADDR 1724
			"00000000000000000000000000000000" , -- ADDR 1725
			"00000000000000000000000000000000" , -- ADDR 1726
			"00000000000000000000000000000000" , -- ADDR 1727
			"00000000000000000000000000000000" , -- ADDR 1728
			"00000000000000000000000000000000" , -- ADDR 1729
			"00000000000000000000000000000000" , -- ADDR 1730
			"00000000000000000000000000000000" , -- ADDR 1731
			"00000000000000000000000000000000" , -- ADDR 1732
			"00000000000000000000000000000000" , -- ADDR 1733
			"00000000000000000000000000000000" , -- ADDR 1734
			"00000000000000000000000000000000" , -- ADDR 1735
			"00000000000000000000000000000000" , -- ADDR 1736
			"00000000000000000000000000000000" , -- ADDR 1737
			"00000000000000000000000000000000" , -- ADDR 1738
			"00000000000000000000000000000000" , -- ADDR 1739
			"00000000000000000000000000000000" , -- ADDR 1740
			"00000000000000000000000000000000" , -- ADDR 1741
			"00000000000000000000000000000000" , -- ADDR 1742
			"00000000000000000000000000000000" , -- ADDR 1743
			"00000000000000000000000000000000" , -- ADDR 1744
			"00000000000000000000000000000000" , -- ADDR 1745
			"00000000000000000000000000000000" , -- ADDR 1746
			"00000000000000000000000000000000" , -- ADDR 1747
			"00000000000000000000000000000000" , -- ADDR 1748
			"00000000000000000000000000000000" , -- ADDR 1749
			"00000000000000000000000000000000" , -- ADDR 1750
			"00000000000000000000000000000000" , -- ADDR 1751
			"00000000000000000000000000000000" , -- ADDR 1752
			"00000000000000000000000000000000" , -- ADDR 1753
			"00000000000000000000000000000000" , -- ADDR 1754
			"00000000000000000000000000000000" , -- ADDR 1755
			"00000000000000000000000000000000" , -- ADDR 1756
			"00000000000000000000000000000000" , -- ADDR 1757
			"00000000000000000000000000000000" , -- ADDR 1758
			"00000000000000000000000000000000" , -- ADDR 1759
			"00000000000000000000000000000000" , -- ADDR 1760
			"00000000000000000000000000000000" , -- ADDR 1761
			"00000000000000000000000000000000" , -- ADDR 1762
			"00000000000000000000000000000000" , -- ADDR 1763
			"00000000000000000000000000000000" , -- ADDR 1764
			"00000000000000000000000000000000" , -- ADDR 1765
			"00000000000000000000000000000000" , -- ADDR 1766
			"00000000000000000000000000000000" , -- ADDR 1767
			"00000000000000000000000000000000" , -- ADDR 1768
			"00000000000000000000000000000000" , -- ADDR 1769
			"00000000000000000000000000000000" , -- ADDR 1770
			"00000000000000000000000000000000" , -- ADDR 1771
			"00000000000000000000000000000000" , -- ADDR 1772
			"00000000000000000000000000000000" , -- ADDR 1773
			"00000000000000000000000000000000" , -- ADDR 1774
			"00000000000000000000000000000000" , -- ADDR 1775
			"00000000000000000000000000000000" , -- ADDR 1776
			"00000000000000000000000000000000" , -- ADDR 1777
			"00000000000000000000000000000000" , -- ADDR 1778
			"00000000000000000000000000000000" , -- ADDR 1779
			"00000000000000000000000000000000" , -- ADDR 1780
			"00000000000000000000000000000000" , -- ADDR 1781
			"00000000000000000000000000000000" , -- ADDR 1782
			"00000000000000000000000000000000" , -- ADDR 1783
			"00000000000000000000000000000000" , -- ADDR 1784
			"00000000000000000000000000000000" , -- ADDR 1785
			"00000000000000000000000000000000" , -- ADDR 1786
			"00000000000000000000000000000000" , -- ADDR 1787
			"00000000000000000000000000000000" , -- ADDR 1788
			"00000000000000000000000000000000" , -- ADDR 1789
			"00000000000000000000000000000000" , -- ADDR 1790
			"00000000000000000000000000000000" , -- ADDR 1791
			"00000000000000000000000000000000" , -- ADDR 1792
			"00000000000000000000000000000000" , -- ADDR 1793
			"00000000000000000000000000000000" , -- ADDR 1794
			"00000000000000000000000000000000" , -- ADDR 1795
			"00000000000000000000000000000000" , -- ADDR 1796
			"00000000000000000000000000000000" , -- ADDR 1797
			"00000000000000000000000000000000" , -- ADDR 1798
			"00000000000000000000000000000000" , -- ADDR 1799
			"00000000000000000000000000000000" , -- ADDR 1800
			"00000000000000000000000000000000" , -- ADDR 1801
			"00000000000000000000000000000000" , -- ADDR 1802
			"00000000000000000000000000000000" , -- ADDR 1803
			"00000000000000000000000000000000" , -- ADDR 1804
			"00000000000000000000000000000000" , -- ADDR 1805
			"00000000000000000000000000000000" , -- ADDR 1806
			"00000000000000000000000000000000" , -- ADDR 1807
			"00000000000000000000000000000000" , -- ADDR 1808
			"00000000000000000000000000000000" , -- ADDR 1809
			"00000000000000000000000000000000" , -- ADDR 1810
			"00000000000000000000000000000000" , -- ADDR 1811
			"00000000000000000000000000000000" , -- ADDR 1812
			"00000000000000000000000000000000" , -- ADDR 1813
			"00000000000000000000000000000000" , -- ADDR 1814
			"00000000000000000000000000000000" , -- ADDR 1815
			"00000000000000000000000000000000" , -- ADDR 1816
			"00000000000000000000000000000000" , -- ADDR 1817
			"00000000000000000000000000000000" , -- ADDR 1818
			"00000000000000000000000000000000" , -- ADDR 1819
			"00000000000000000000000000000000" , -- ADDR 1820
			"00000000000000000000000000000000" , -- ADDR 1821
			"00000000000000000000000000000000" , -- ADDR 1822
			"00000000000000000000000000000000" , -- ADDR 1823
			"00000000000000000000000000000000" , -- ADDR 1824
			"00000000000000000000000000000000" , -- ADDR 1825
			"00000000000000000000000000000000" , -- ADDR 1826
			"00000000000000000000000000000000" , -- ADDR 1827
			"00000000000000000000000000000000" , -- ADDR 1828
			"00000000000000000000000000000000" , -- ADDR 1829
			"00000000000000000000000000000000" , -- ADDR 1830
			"00000000000000000000000000000000" , -- ADDR 1831
			"00000000000000000000000000000000" , -- ADDR 1832
			"00000000000000000000000000000000" , -- ADDR 1833
			"00000000000000000000000000000000" , -- ADDR 1834
			"00000000000000000000000000000000" , -- ADDR 1835
			"00000000000000000000000000000000" , -- ADDR 1836
			"00000000000000000000000000000000" , -- ADDR 1837
			"00000000000000000000000000000000" , -- ADDR 1838
			"00000000000000000000000000000000" , -- ADDR 1839
			"00000000000000000000000000000000" , -- ADDR 1840
			"00000000000000000000000000000000" , -- ADDR 1841
			"00000000000000000000000000000000" , -- ADDR 1842
			"00000000000000000000000000000000" , -- ADDR 1843
			"00000000000000000000000000000000" , -- ADDR 1844
			"00000000000000000000000000000000" , -- ADDR 1845
			"00000000000000000000000000000000" , -- ADDR 1846
			"00000000000000000000000000000000" , -- ADDR 1847
			"00000000000000000000000000000000" , -- ADDR 1848
			"00000000000000000000000000000000" , -- ADDR 1849
			"00000000000000000000000000000000" , -- ADDR 1850
			"00000000000000000000000000000000" , -- ADDR 1851
			"00000000000000000000000000000000" , -- ADDR 1852
			"00000000000000000000000000000000" , -- ADDR 1853
			"00000000000000000000000000000000" , -- ADDR 1854
			"00000000000000000000000000000000" , -- ADDR 1855
			"00000000000000000000000000000000" , -- ADDR 1856
			"00000000000000000000000000000000" , -- ADDR 1857
			"00000000000000000000000000000000" , -- ADDR 1858
			"00000000000000000000000000000000" , -- ADDR 1859
			"00000000000000000000000000000000" , -- ADDR 1860
			"00000000000000000000000000000000" , -- ADDR 1861
			"00000000000000000000000000000000" , -- ADDR 1862
			"00000000000000000000000000000000" , -- ADDR 1863
			"00000000000000000000000000000000" , -- ADDR 1864
			"00000000000000000000000000000000" , -- ADDR 1865
			"00000000000000000000000000000000" , -- ADDR 1866
			"00000000000000000000000000000000" , -- ADDR 1867
			"00000000000000000000000000000000" , -- ADDR 1868
			"00000000000000000000000000000000" , -- ADDR 1869
			"00000000000000000000000000000000" , -- ADDR 1870
			"00000000000000000000000000000000" , -- ADDR 1871
			"00000000000000000000000000000000" , -- ADDR 1872
			"00000000000000000000000000000000" , -- ADDR 1873
			"00000000000000000000000000000000" , -- ADDR 1874
			"00000000000000000000000000000000" , -- ADDR 1875
			"00000000000000000000000000000000" , -- ADDR 1876
			"00000000000000000000000000000000" , -- ADDR 1877
			"00000000000000000000000000000000" , -- ADDR 1878
			"00000000000000000000000000000000" , -- ADDR 1879
			"00000000000000000000000000000000" , -- ADDR 1880
			"00000000000000000000000000000000" , -- ADDR 1881
			"00000000000000000000000000000000" , -- ADDR 1882
			"00000000000000000000000000000000" , -- ADDR 1883
			"00000000000000000000000000000000" , -- ADDR 1884
			"00000000000000000000000000000000" , -- ADDR 1885
			"00000000000000000000000000000000" , -- ADDR 1886
			"00000000000000000000000000000000" , -- ADDR 1887
			"00000000000000000000000000000000" , -- ADDR 1888
			"00000000000000000000000000000000" , -- ADDR 1889
			"00000000000000000000000000000000" , -- ADDR 1890
			"00000000000000000000000000000000" , -- ADDR 1891
			"00000000000000000000000000000000" , -- ADDR 1892
			"00000000000000000000000000000000" , -- ADDR 1893
			"00000000000000000000000000000000" , -- ADDR 1894
			"00000000000000000000000000000000" , -- ADDR 1895
			"00000000000000000000000000000000" , -- ADDR 1896
			"00000000000000000000000000000000" , -- ADDR 1897
			"00000000000000000000000000000000" , -- ADDR 1898
			"00000000000000000000000000000000" , -- ADDR 1899
			"00000000000000000000000000000000" , -- ADDR 1900
			"00000000000000000000000000000000" , -- ADDR 1901
			"00000000000000000000000000000000" , -- ADDR 1902
			"00000000000000000000000000000000" , -- ADDR 1903
			"00000000000000000000000000000000" , -- ADDR 1904
			"00000000000000000000000000000000" , -- ADDR 1905
			"00000000000000000000000000000000" , -- ADDR 1906
			"00000000000000000000000000000000" , -- ADDR 1907
			"00000000000000000000000000000000" , -- ADDR 1908
			"00000000000000000000000000000000" , -- ADDR 1909
			"00000000000000000000000000000000" , -- ADDR 1910
			"00000000000000000000000000000000" , -- ADDR 1911
			"00000000000000000000000000000000" , -- ADDR 1912
			"00000000000000000000000000000000" , -- ADDR 1913
			"00000000000000000000000000000000" , -- ADDR 1914
			"00000000000000000000000000000000" , -- ADDR 1915
			"00000000000000000000000000000000" , -- ADDR 1916
			"00000000000000000000000000000000" , -- ADDR 1917
			"00000000000000000000000000000000" , -- ADDR 1918
			"00000000000000000000000000000000" , -- ADDR 1919
			"00000000000000000000000000000000" , -- ADDR 1920
			"00000000000000000000000000000000" , -- ADDR 1921
			"00000000000000000000000000000000" , -- ADDR 1922
			"00000000000000000000000000000000" , -- ADDR 1923
			"00000000000000000000000000000000" , -- ADDR 1924
			"00000000000000000000000000000000" , -- ADDR 1925
			"00000000000000000000000000000000" , -- ADDR 1926
			"00000000000000000000000000000000" , -- ADDR 1927
			"00000000000000000000000000000000" , -- ADDR 1928
			"00000000000000000000000000000000" , -- ADDR 1929
			"00000000000000000000000000000000" , -- ADDR 1930
			"00000000000000000000000000000000" , -- ADDR 1931
			"00000000000000000000000000000000" , -- ADDR 1932
			"00000000000000000000000000000000" , -- ADDR 1933
			"00000000000000000000000000000000" , -- ADDR 1934
			"00000000000000000000000000000000" , -- ADDR 1935
			"00000000000000000000000000000000" , -- ADDR 1936
			"00000000000000000000000000000000" , -- ADDR 1937
			"00000000000000000000000000000000" , -- ADDR 1938
			"00000000000000000000000000000000" , -- ADDR 1939
			"00000000000000000000000000000000" , -- ADDR 1940
			"00000000000000000000000000000000" , -- ADDR 1941
			"00000000000000000000000000000000" , -- ADDR 1942
			"00000000000000000000000000000000" , -- ADDR 1943
			"00000000000000000000000000000000" , -- ADDR 1944
			"00000000000000000000000000000000" , -- ADDR 1945
			"00000000000000000000000000000000" , -- ADDR 1946
			"00000000000000000000000000000000" , -- ADDR 1947
			"00000000000000000000000000000000" , -- ADDR 1948
			"00000000000000000000000000000000" , -- ADDR 1949
			"00000000000000000000000000000000" , -- ADDR 1950
			"00000000000000000000000000000000" , -- ADDR 1951
			"00000000000000000000000000000000" , -- ADDR 1952
			"00000000000000000000000000000000" , -- ADDR 1953
			"00000000000000000000000000000000" , -- ADDR 1954
			"00000000000000000000000000000000" , -- ADDR 1955
			"00000000000000000000000000000000" , -- ADDR 1956
			"00000000000000000000000000000000" , -- ADDR 1957
			"00000000000000000000000000000000" , -- ADDR 1958
			"00000000000000000000000000000000" , -- ADDR 1959
			"00000000000000000000000000000000" , -- ADDR 1960
			"00000000000000000000000000000000" , -- ADDR 1961
			"00000000000000000000000000000000" , -- ADDR 1962
			"00000000000000000000000000000000" , -- ADDR 1963
			"00000000000000000000000000000000" , -- ADDR 1964
			"00000000000000000000000000000000" , -- ADDR 1965
			"00000000000000000000000000000000" , -- ADDR 1966
			"00000000000000000000000000000000" , -- ADDR 1967
			"00000000000000000000000000000000" , -- ADDR 1968
			"00000000000000000000000000000000" , -- ADDR 1969
			"00000000000000000000000000000000" , -- ADDR 1970
			"00000000000000000000000000000000" , -- ADDR 1971
			"00000000000000000000000000000000" , -- ADDR 1972
			"00000000000000000000000000000000" , -- ADDR 1973
			"00000000000000000000000000000000" , -- ADDR 1974
			"00000000000000000000000000000000" , -- ADDR 1975
			"00000000000000000000000000000000" , -- ADDR 1976
			"00000000000000000000000000000000" , -- ADDR 1977
			"00000000000000000000000000000000" , -- ADDR 1978
			"00000000000000000000000000000000" , -- ADDR 1979
			"00000000000000000000000000000000" , -- ADDR 1980
			"00000000000000000000000000000000" , -- ADDR 1981
			"00000000000000000000000000000000" , -- ADDR 1982
			"00000000000000000000000000000000" , -- ADDR 1983
			"00000000000000000000000000000000" , -- ADDR 1984
			"00000000000000000000000000000000" , -- ADDR 1985
			"00000000000000000000000000000000" , -- ADDR 1986
			"00000000000000000000000000000000" , -- ADDR 1987
			"00000000000000000000000000000000" , -- ADDR 1988
			"00000000000000000000000000000000" , -- ADDR 1989
			"00000000000000000000000000000000" , -- ADDR 1990
			"00000000000000000000000000000000" , -- ADDR 1991
			"00000000000000000000000000000000" , -- ADDR 1992
			"00000000000000000000000000000000" , -- ADDR 1993
			"00000000000000000000000000000000" , -- ADDR 1994
			"00000000000000000000000000000000" , -- ADDR 1995
			"00000000000000000000000000000000" , -- ADDR 1996
			"00000000000000000000000000000000" , -- ADDR 1997
			"00000000000000000000000000000000" , -- ADDR 1998
			"00000000000000000000000000000000" , -- ADDR 1999
			"00000000000000000000000000000000" , -- ADDR 2000
			"00000000000000000000000000000000" , -- ADDR 2001
			"00000000000000000000000000000000" , -- ADDR 2002
			"00000000000000000000000000000000" , -- ADDR 2003
			"00000000000000000000000000000000" , -- ADDR 2004
			"00000000000000000000000000000000" , -- ADDR 2005
			"00000000000000000000000000000000" , -- ADDR 2006
			"00000000000000000000000000000000" , -- ADDR 2007
			"00000000000000000000000000000000" , -- ADDR 2008
			"00000000000000000000000000000000" , -- ADDR 2009
			"00000000000000000000000000000000" , -- ADDR 2010
			"00000000000000000000000000000000" , -- ADDR 2011
			"00000000000000000000000000000000" , -- ADDR 2012
			"00000000000000000000000000000000" , -- ADDR 2013
			"00000000000000000000000000000000" , -- ADDR 2014
			"00000000000000000000000000000000" , -- ADDR 2015
			"00000000000000000000000000000000" , -- ADDR 2016
			"00000000000000000000000000000000" , -- ADDR 2017
			"00000000000000000000000000000000" , -- ADDR 2018
			"00000000000000000000000000000000" , -- ADDR 2019
			"00000000000000000000000000000000" , -- ADDR 2020
			"00000000000000000000000000000000" , -- ADDR 2021
			"00000000000000000000000000000000" , -- ADDR 2022
			"00000000000000000000000000000000" , -- ADDR 2023
			"00000000000000000000000000000000" , -- ADDR 2024
			"00000000000000000000000000000000" , -- ADDR 2025
			"00000000000000000000000000000000" , -- ADDR 2026
			"00000000000000000000000000000000" , -- ADDR 2027
			"00000000000000000000000000000000" , -- ADDR 2028
			"00000000000000000000000000000000" , -- ADDR 2029
			"00000000000000000000000000000000" , -- ADDR 2030
			"00000000000000000000000000000000" , -- ADDR 2031
			"00000000000000000000000000000000" , -- ADDR 2032
			"00000000000000000000000000000000" , -- ADDR 2033
			"00000000000000000000000000000000" , -- ADDR 2034
			"00000000000000000000000000000000" , -- ADDR 2035
			"00000000000000000000000000000000" , -- ADDR 2036
			"00000000000000000000000000000000" , -- ADDR 2037
			"00000000000000000000000000000000" , -- ADDR 2038
			"00000000000000000000000000000000" , -- ADDR 2039
			"00000000000000000000000000000000" , -- ADDR 2040
			"00000000000000000000000000000000" , -- ADDR 2041
			"00000000000000000000000000000000" , -- ADDR 2042
			"00000000000000000000000000000000" , -- ADDR 2043
			"00000000000000000000000000000000" , -- ADDR 2044
			"00000000000000000000000000000000" , -- ADDR 2045
			"00000000000000000000000000000000" , -- ADDR 2046
			"00000000000000000000000000000000"   -- ADDR 2047
			);
			
begin
	
	process (CLK)
	begin
		if (rising_edge(CLK)) then
			-- In the case of Altera Quartus, it is extremely essential that the output assignment stays in the process.
			-- Otherwise, Altera Quartus will not infer the VHDL code as ROM.
			-- However, in the case of Xilinx ISE, it does not matter whether the output assignment stays in the process
			-- or outside of it with synchronization to the clock pulse by another signal. The VHDL code will infer as ROM anyway.
			DATA <= ROM (to_integer(unsigned(ADDR)));
		end if;
	end process;
	
end Behavioral;

-- Extremely important: In order for Altera Quartus to infer the VHDL code as ROM, the setting in the path
-- "Assignments/Device�/Device and Pin Options�/Configuration/Configuration mode" must be changed to
-- "Single Uncompressed Image with memory initialization (512 Kbits UFM)".