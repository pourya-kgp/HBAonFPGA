----------------------------------------------------------------------------------------------------
-- Author           : Pourya Khodagholipour (P.KH)
-- Project Name     : HBA (Hardware Bee Algorithm)
-- File Name        : TSP_Dist_One_Port_ROM_Sync
-- Module Name      : TSP_Dist_One_Port_ROM_Sync
-- HDL Standard     : VHDL
-- Approach         : Behavioral
-- Description      : Single-port ROM with synchronous read (Block RAM)
-- Comments         : st70 Database Distance matrix
-- Dependencies     : ---
-- Target Devices   : Virtex 5 - XC5VLX330
-- Speed Estimation : ---
-- Area  Estimation : 4 RAM/FIFO
-- Tools            : ISE Design Suite v14.7 - Altera Quartus 16.1 Lite
-- Module Version   : 
-- Creation Date    : 2016/08
-- Revision Date    : 2024/07/08
----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity TSP_Dist_One_Port_ROM_Sync is
	generic (
				ADDR_WIDTH : natural := 12;
				DATA_WIDTH : natural := 32);
	port    (
				CLK        : in  std_logic;
				ADDR       : in  std_logic_vector (ADDR_WIDTH-1 downto 0);
				DATA       : out std_logic_vector (DATA_WIDTH-1 downto 0));
end TSP_Dist_One_Port_ROM_Sync;

architecture Behavioral of TSP_Dist_One_Port_ROM_Sync is

	type ROM_Type is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector (DATA_WIDTH-1 downto 0);
	constant ROM : ROM_Type := (
			"11111111111111111111111111111111" , -- ADDR 0
			"00000000000000001110011101000011" , -- ADDR 1
			"00000000000000010001110111010011" , -- ADDR 2
			"00000000000000001101010100111101" , -- ADDR 3
			"00000000000000001000000101100001" , -- ADDR 4
			"00000000000000001101000001011011" , -- ADDR 5
			"00000000000000001111101100100000" , -- ADDR 6
			"00000000000000010011101000011011" , -- ADDR 7
			"00000000000000010011101010010001" , -- ADDR 8
			"00000000000000001000111000110001" , -- ADDR 9
			"00000000000000001110101111110111" , -- ADDR 10
			"00000000000000001101111010110001" , -- ADDR 11
			"00000000000000000011100011100000" , -- ADDR 12
			"00000000000000010101011111000000" , -- ADDR 13
			"00000000000000001100001010011100" , -- ADDR 14
			"00000000000000000010000110011010" , -- ADDR 15
			"00000000000000010000000000010000" , -- ADDR 16
			"00000000000000001101101101001111" , -- ADDR 17
			"00000000000000010000100110111101" , -- ADDR 18
			"00000000000000010111001100101101" , -- ADDR 19
			"00000000000000001111101001000110" , -- ADDR 20
			"00000000000000000110010101010110" , -- ADDR 21
			"00000000000000000010000101100000" , -- ADDR 22
			"00000000000000001100011101011111" , -- ADDR 23
			"00000000000000011001101110110010" , -- ADDR 24
			"00000000000000010011110110101000" , -- ADDR 25
			"00000000000000010110110011100000" , -- ADDR 26
			"00000000000000010100100000101100" , -- ADDR 27
			"00000000000000000011011100111110" , -- ADDR 28
			"00000000000000010110110011111010" , -- ADDR 29
			"00000000000000000100110011110010" , -- ADDR 30
			"00000000000000010000101111110001" , -- ADDR 31
			"00000000000000001110101011101101" , -- ADDR 32
			"00000000000000001111110001111101" , -- ADDR 33
			"00000000000000000111111100111101" , -- ADDR 34
			"00000000000000000001000010010011" , -- ADDR 35
			"00000000000000000101000010001000" , -- ADDR 36
			"00000000000000000100100010101001" , -- ADDR 37
			"00000000000000010111001111101010" , -- ADDR 38
			"00000000000000010101110111010010" , -- ADDR 39
			"00000000000000001110010111101000" , -- ADDR 40
			"00000000000000001110101001101000" , -- ADDR 41
			"00000000000000010000001000110010" , -- ADDR 42
			"00000000000000010011010001000110" , -- ADDR 43
			"00000000000000010111111010011000" , -- ADDR 44
			"00000000000000011000001010111101" , -- ADDR 45
			"00000000000000000011000011110010" , -- ADDR 46
			"00000000000000010000000011001110" , -- ADDR 47
			"00000000000000010110001010110010" , -- ADDR 48
			"00000000000000000111011100010000" , -- ADDR 49
			"00000000000000001010101100110101" , -- ADDR 50
			"00000000000000001010001110001101" , -- ADDR 51
			"00000000000000001000010010100100" , -- ADDR 52
			"00000000000000010000100011011001" , -- ADDR 53
			"00000000000000010111010000101001" , -- ADDR 54
			"00000000000000001100111001000010" , -- ADDR 55
			"00000000000000001010101100110101" , -- ADDR 56
			"00000000000000000101001100001100" , -- ADDR 57
			"00000000000000000110011010001001" , -- ADDR 58
			"00000000000000001100010000100010" , -- ADDR 59
			"00000000000000010101011001110000" , -- ADDR 60
			"00000000000000010011000010100011" , -- ADDR 61
			"00000000000000000111010101000001" , -- ADDR 62
			"00000000000000001101011101101001" , -- ADDR 63
			"00000000000000001011111110010001" , -- ADDR 64
			"00000000000000000111011111010100" , -- ADDR 65
			"00000000000000001110110110011100" , -- ADDR 66
			"00000000000000010011001100110101" , -- ADDR 67
			"00000000000000000101001111011111" , -- ADDR 68
			"00000000000000000100111010000100" , -- ADDR 69
			"00000000000000000100101111011000" , -- ADDR 70
			"00000000000000000010000101100000" , -- ADDR 71
			"00000000000000001010011000011001" , -- ADDR 72
			"00000000000000000101011101011001" , -- ADDR 73
			"00000000000000000001001111101011" , -- ADDR 74
			"00000000000000000101011000000111" , -- ADDR 75
			"00000000000000001100110100010010" , -- ADDR 76
			"00000000000000001011100001100010" , -- ADDR 77
			"00000000000000010011111110110001" , -- ADDR 78
			"00000000000000001100110010101001" , -- ADDR 79
			"00000000000000001100111100101110" , -- ADDR 80
			"00000000000000001000100001000110" , -- ADDR 81
			"00000000000000000101101110000111" , -- ADDR 82
			"00000000000000001101111000011011" , -- ADDR 83
			"00000000000000001001110100001000" , -- ADDR 84
			"00000000000000000010111100001010" , -- ADDR 85
			"00000000000000000011001011001000" , -- ADDR 86
			"00000000000000001010010001000000" , -- ADDR 87
			"00000000000000001100101110111010" , -- ADDR 88
			"00000000000000001000010110111010" , -- ADDR 89
			"00000000000000001100011000000111" , -- ADDR 90
			"00000000000000000100110110001001" , -- ADDR 91
			"00000000000000010011100101100111" , -- ADDR 92
			"00000000000000000101011001111000" , -- ADDR 93
			"00000000000000001110001111000110" , -- ADDR 94
			"00000000000000000110011000111101" , -- ADDR 95
			"00000000000000001101011011111100" , -- ADDR 96
			"00000000000000001010101100110101" , -- ADDR 97
			"00000000000000001011111110010001" , -- ADDR 98
			"00000000000000000011001011101110" , -- ADDR 99
			"00000000000000001111001010010001" , -- ADDR 100
			"00000000000000001100111110011111" , -- ADDR 101
			"00000000000000001100000010111000" , -- ADDR 102
			"00000000000000001110111111010000" , -- ADDR 103
			"00000000000000001101010010000110" , -- ADDR 104
			"00000000000000001010010100111001" , -- ADDR 105
			"00000000000000010010001111100110" , -- ADDR 106
			"00000000000000001111100001010001" , -- ADDR 107
			"00000000000000000110010110100011" , -- ADDR 108
			"00000000000000000100001101101111" , -- ADDR 109
			"00000000000000001000111010010001" , -- ADDR 110
			"00000000000000001000100010111000" , -- ADDR 111
			"00000000000000010001110001100001" , -- ADDR 112
			"00000000000000001111110010010101" , -- ADDR 113
			"00000000000000001100011100101110" , -- ADDR 114
			"00000000000000010011100010111000" , -- ADDR 115
			"00000000000000000111101110000111" , -- ADDR 116
			"00000000000000001101000111111111" , -- ADDR 117
			"00000000000000010000001011101111" , -- ADDR 118
			"00000000000000001100001001001011" , -- ADDR 119
			"00000000000000001000010010010101" , -- ADDR 120
			"00000000000000010001100001111101" , -- ADDR 121
			"00000000000000001000111101101011" , -- ADDR 122
			"00000000000000010001110011110001" , -- ADDR 123
			"00000000000000000101100100111111" , -- ADDR 124
			"00000000000000001101000101100000" , -- ADDR 125
			"00000000000000001001000010010110" , -- ADDR 126
			"00000000000000001101011101110010" , -- ADDR 127
			"00000000000000001111111011100101" , -- ADDR 128
			"00000000000000010010010111101000" , -- ADDR 129
			"00000000000000000111100100101000" , -- ADDR 130
			"00000000000000010110110110100110" , -- ADDR 131
			"00000000000000010010100111110100" , -- ADDR 132
			"00000000000000000110111111011100" , -- ADDR 133
			"00000000000000010010011111111001" , -- ADDR 134
			"00000000000000001001001101101000" , -- ADDR 135
			"00000000000000001011011111111000" , -- ADDR 136
			"00000000000000001101011101101001" , -- ADDR 137
			"00000000000000000100101100100011" , -- ADDR 138
			"00000000000000001011111001110010" , -- ADDR 139
			"00000000000000000101100100101001" , -- ADDR 140
			"00000000000000000011111110010111" , -- ADDR 141
			"00000000000000000010110110001110" , -- ADDR 142
			"00000000000000001001100001011000" , -- ADDR 143
			"00000000000000001100100110101000" , -- ADDR 144
			"00000000000000010011111010011110" , -- ADDR 145
			"00000000000000001011111010111010" , -- ADDR 146
			"00000000000000010000111111010000" , -- ADDR 147
			"00000000000000000011110111000011" , -- ADDR 148
			"00000000000000001010011100110010" , -- ADDR 149
			"00000000000000010000110110111011" , -- ADDR 150
			"00000000000000000111101010011001" , -- ADDR 151
			"00000000000000000100001010000101" , -- ADDR 152
			"00000000000000000110001110010111" , -- ADDR 153
			"00000000000000000101101000101111" , -- ADDR 154
			"00000000000000001011001000110010" , -- ADDR 155
			"00000000000000001100010100111000" , -- ADDR 156
			"00000000000000001111111000000111" , -- ADDR 157
			"00000000000000001001100100100101" , -- ADDR 158
			"00000000000000001111110011111001" , -- ADDR 159
			"00000000000000000100100011111010" , -- ADDR 160
			"00000000000000001010000111011101" , -- ADDR 161
			"00000000000000000011001000000110" , -- ADDR 162
			"00000000000000010001011110010000" , -- ADDR 163
			"00000000000000000101111101011101" , -- ADDR 164
			"00000000000000010000001011101111" , -- ADDR 165
			"00000000000000000001100100000011" , -- ADDR 166
			"00000000000000001110010010011011" , -- ADDR 167
			"00000000000000001011010110110111" , -- ADDR 168
			"00000000000000010000101000111010" , -- ADDR 169
			"00000000000000010010100011111010" , -- ADDR 170
			"00000000000000001111100001010001" , -- ADDR 171
			"00000000000000001110001111000110" , -- ADDR 172
			"00000000000000001110111011001011" , -- ADDR 173
			"00000000000000001100000001100110" , -- ADDR 174
			"00000000000000000101001011011101" , -- ADDR 175
			"00000000000000000011011111101110" , -- ADDR 176
			"00000000000000000110100100101110" , -- ADDR 177
			"00000000000000000100010100111000" , -- ADDR 178
			"00000000000000001110001000001111" , -- ADDR 179
			"00000000000000001011100110110011" , -- ADDR 180
			"00000000000000001111010111111000" , -- ADDR 181
			"00000000000000010010111101100010" , -- ADDR 182
			"00000000000000000110001010010111" , -- ADDR 183
			"00000000000000001110101000100110" , -- ADDR 184
			"00000000000000010000110100010100" , -- ADDR 185
			"00000000000000001100101100101010" , -- ADDR 186
			"00000000000000001010010001001011" , -- ADDR 187
			"00000000000000010000011000101111" , -- ADDR 188
			"00000000000000001000000101100001" , -- ADDR 189
			"00000000000000010001111101010001" , -- ADDR 190
			"00000000000000001010010001001011" , -- ADDR 191
			"00000000000000001111010010100010" , -- ADDR 192
			"00000000000000001101010001000110" , -- ADDR 193
			"00000000000000001101010011011001" , -- ADDR 194
			"00000000000000001100101100101010" , -- ADDR 195
			"00000000000000010000100001011100" , -- ADDR 196
			"00000000000000001011101110110100" , -- ADDR 197
			"00000000000000010111110101010001" , -- ADDR 198
			"00000000000000010011001100110101" , -- ADDR 199
			"00000000000000001010110011111011" , -- ADDR 200
			"00000000000000010010000111011010" , -- ADDR 201
			"00000000000000000101001110000010" , -- ADDR 202
			"00000000000000001111110000011001" , -- ADDR 203
			"00000000000000010001101101110111" , -- ADDR 204
			"00000000000000001000011101011111" , -- ADDR 205
			"00000000000000000011011011010100" , -- ADDR 206
			"00000000000000000010111100001010" , -- ADDR 207
			"00000000000000000110010101101010" , -- ADDR 208
			"00000000000000001011010000010010" , -- ADDR 209
			"00000000000000001001100010001011" , -- ADDR 210
			"00000000000000010001111010001011" , -- ADDR 211
			"00000000000000001010101110011100" , -- ADDR 212
			"00000000000000001100010010110111" , -- ADDR 213
			"00000000000000001000100001110000" , -- ADDR 214
			"00000000000000000110101101000011" , -- ADDR 215
			"00000000000000001100100000101101" , -- ADDR 216
			"00000000000000000111111111110101" , -- ADDR 217
			"00000000000000000001000101111000" , -- ADDR 218
			"00000000000000000101010000100101" , -- ADDR 219
			"00000000000000001010010011011010" , -- ADDR 220
			"00000000000000001010101111101011" , -- ADDR 221
			"00000000000000000111101000011001" , -- ADDR 222
			"00000000000000001011010010111111" , -- ADDR 223
			"00000000000000000101111001111011" , -- ADDR 224
			"00000000000000010010001000000011" , -- ADDR 225
			"00000000000000000110111010001110" , -- ADDR 226
			"00000000000000001101000010100101" , -- ADDR 227
			"00000000000000000111001011110100" , -- ADDR 228
			"00000000000000001100110001111001" , -- ADDR 229
			"00000000000000001010011000110000" , -- ADDR 230
			"00000000000000001011011111100010" , -- ADDR 231
			"00000000000000000011011011010100" , -- ADDR 232
			"00000000000000001101000101100000" , -- ADDR 233
			"00000000000000001010111111010011" , -- ADDR 234
			"00000000000000001100000111110001" , -- ADDR 235
			"00000000000000001101111110000011" , -- ADDR 236
			"00000000000000001011100110010100" , -- ADDR 237
			"00000000000000001001100011001011" , -- ADDR 238
			"00000000000000010000100110100111" , -- ADDR 239
			"00000000000000001101111110110111" , -- ADDR 240
			"00000000000000000100100000000111" , -- ADDR 241
			"00000000000000000010101001000001" , -- ADDR 242
			"00000000000000000111001011100011" , -- ADDR 243
			"00000000000000000111101000001001" , -- ADDR 244
			"00000000000000010000010001010001" , -- ADDR 245
			"00000000000000001110100110101000" , -- ADDR 246
			"00000000000000001011000010100110" , -- ADDR 247
			"00000000000000010001011101011000" , -- ADDR 248
			"00000000000000001001001011010110" , -- ADDR 249
			"00000000000000001011001110111011" , -- ADDR 250
			"00000000000000001110001010011001" , -- ADDR 251
			"00000000000000001010000101111100" , -- ADDR 252
			"00000000000000000110011100100001" , -- ADDR 253
			"00000000000000001111011101110100" , -- ADDR 254
			"00000000000000001010101001010000" , -- ADDR 255
			"00000000000000001111101111110010" , -- ADDR 256
			"00000000000000000110000010110111" , -- ADDR 257
			"00000000000000001011011000111000" , -- ADDR 258
			"00000000000000001000100101100011" , -- ADDR 259
			"00000000000000001011011000010111" , -- ADDR 260
			"00000000000000001110010010011011" , -- ADDR 261
			"00000000000000010000010111111011" , -- ADDR 262
			"00000000000000000111000010111110" , -- ADDR 263
			"00000000000000010100111010000001" , -- ADDR 264
			"00000000000000010000100110100111" , -- ADDR 265
			"00000000000000000110000111111000" , -- ADDR 266
			"00000000000000010000011010011111" , -- ADDR 267
			"00000000000000001000000111011010" , -- ADDR 268
			"00000000000000001011000100101010" , -- ADDR 269
			"00000000000000001101000001110111" , -- ADDR 270
			"00000000000000000110010110010000" , -- ADDR 271
			"00000000000000001011011001001101" , -- ADDR 272
			"00000000000000001110010111001110" , -- ADDR 273
			"00000000000000001011100110110011" , -- ADDR 274
			"00000000000000000001011101110000" , -- ADDR 275
			"00000000000000001010001111111000" , -- ADDR 276
			"00000000000000000110000100000111" , -- ADDR 277
			"00000000000000001001100010001011" , -- ADDR 278
			"00000000000000001110111011001011" , -- ADDR 279
			"00000000000000001011101110110100" , -- ADDR 280
			"00000000000000000110010000100000" , -- ADDR 281
			"00000000000000001000000011011001" , -- ADDR 282
			"00000000000000001000001101000001" , -- ADDR 283
			"00000000000000001101011011011000" , -- ADDR 284
			"00000000000000010000011110001101" , -- ADDR 285
			"00000000000000000111101000001001" , -- ADDR 286
			"00000000000000000110111111011100" , -- ADDR 287
			"00000000000000000110111010100000" , -- ADDR 288
			"00000000000000001011011011111000" , -- ADDR 289
			"00000000000000010001101011100110" , -- ADDR 290
			"00000000000000001111010010100010" , -- ADDR 291
			"00000000000000001110110100111001" , -- ADDR 292
			"00000000000000001110111101101110" , -- ADDR 293
			"00000000000000001001110110101001" , -- ADDR 294
			"00000000000000001111101101111110" , -- ADDR 295
			"00000000000000001001110000011010" , -- ADDR 296
			"00000000000000001011010011110101" , -- ADDR 297
			"00000000000000000111011011111111" , -- ADDR 298
			"00000000000000000111110010010010" , -- ADDR 299
			"00000000000000001100011000000111" , -- ADDR 300
			"00000000000000001001000101100000" , -- ADDR 301
			"00000000000000000011111010000000" , -- ADDR 302
			"00000000000000000111011011001110" , -- ADDR 303
			"00000000000000001111010000010010" , -- ADDR 304
			"00000000000000001101110001110100" , -- ADDR 305
			"00000000000000000111001110101110" , -- ADDR 306
			"00000000000000001000011010000110" , -- ADDR 307
			"00000000000000001000010110111010" , -- ADDR 308
			"00000000000000001100000000001011" , -- ADDR 309
			"00000000000000001111110110000100" , -- ADDR 310
			"00000000000000010000001001010001" , -- ADDR 311
			"00000000000000000101000001101111" , -- ADDR 312
			"00000000000000001010011111111000" , -- ADDR 313
			"00000000000000010001011110111010" , -- ADDR 314
			"00000000000000000010110010001010" , -- ADDR 315
			"00000000000000000110000001111010" , -- ADDR 316
			"00000000000000000010110010001010" , -- ADDR 317
			"00000000000000000010001011110000" , -- ADDR 318
			"00000000000000001001101110101010" , -- ADDR 319
			"00000000000000010011000100010110" , -- ADDR 320
			"00000000000000000111111111110101" , -- ADDR 321
			"00000000000000001010001001111001" , -- ADDR 322
			"00000000000000000011101010011000" , -- ADDR 323
			"00000000000000001000010110011101" , -- ADDR 324
			"00000000000000000100111100011000" , -- ADDR 325
			"00000000000000001101010101110100" , -- ADDR 326
			"00000000000000001011110010101101" , -- ADDR 327
			"00000000000000000111100110101001" , -- ADDR 328
			"00000000000000001100011110010000" , -- ADDR 329
			"00000000000000001000011010000110" , -- ADDR 330
			"00000000000000000110010110010000" , -- ADDR 331
			"00000000000000001001010001111101" , -- ADDR 332
			"00000000000000001011101110000000" , -- ADDR 333
			"00000000000000001001101110010001" , -- ADDR 334
			"00000000000000001010111111001000" , -- ADDR 335
			"00000000000000000110000001111010" , -- ADDR 336
			"00000000000000001000001010001110" , -- ADDR 337
			"00000000000000001000011001101001" , -- ADDR 338
			"00000000000000000111000010101100" , -- ADDR 339
			"00000000000000001110110101001001" , -- ADDR 340
			"00000000000000000111010110000011" , -- ADDR 341
			"00000000000000001100111010111100" , -- ADDR 342
			"00000000000000001000101010110111" , -- ADDR 343
			"00000000000000001001101010001000" , -- ADDR 344
			"00000000000000001011101110001010" , -- ADDR 345
			"00000000000000000100110011110010" , -- ADDR 346
			"00000000000000000010100011001000" , -- ADDR 347
			"00000000000000001000100101100011" , -- ADDR 348
			"00000000000000001010010011001110" , -- ADDR 349
			"00000000000000000111010100110000" , -- ADDR 350
			"00000000000000001000100010101010" , -- ADDR 351
			"00000000000000001011001101000011" , -- ADDR 352
			"00000000000000001000111101010000" , -- ADDR 353
			"00000000000000001111010011011010" , -- ADDR 354
			"00000000000000001001010110010000" , -- ADDR 355
			"00000000000000001010110000001101" , -- ADDR 356
			"00000000000000001000101010110111" , -- ADDR 357
			"00000000000000001101010111111101" , -- ADDR 358
			"00000000000000001001110010110000" , -- ADDR 359
			"00000000000000001100011100111000" , -- ADDR 360
			"00000000000000000101001011011101" , -- ADDR 361
			"00000000000000001001101110101010" , -- ADDR 362
			"00000000000000000111100100011000" , -- ADDR 363
			"00000000000000001101110110010111" , -- ADDR 364
			"00000000000000001101110110001111" , -- ADDR 365
			"00000000000000001010000100001111" , -- ADDR 366
			"00000000000000001010001010011101" , -- ADDR 367
			"00000000000000001101100010100110" , -- ADDR 368
			"00000000000000001011000110101110" , -- ADDR 369
			"00000000000000000001100100000011" , -- ADDR 370
			"00000000000000000010000110011010" , -- ADDR 371
			"00000000000000000100001100110101" , -- ADDR 372
			"00000000000000000110010001101110" , -- ADDR 373
			"00000000000000001101011010000110" , -- ADDR 374
			"00000000000000001100010010011001" , -- ADDR 375
			"00000000000000001010010000010000" , -- ADDR 376
			"00000000000000001110001101000101" , -- ADDR 377
			"00000000000000001011011001100010" , -- ADDR 378
			"00000000000000001001000100000001" , -- ADDR 379
			"00000000000000001011011001001101" , -- ADDR 380
			"00000000000000000111010000000010" , -- ADDR 381
			"00000000000000000100111010000100" , -- ADDR 382
			"00000000000000001100000101000101" , -- ADDR 383
			"00000000000000001101001000110110" , -- ADDR 384
			"00000000000000001100101111101010" , -- ADDR 385
			"00000000000000001000101000011011" , -- ADDR 386
			"00000000000000001001110101000110" , -- ADDR 387
			"00000000000000001001110100100000" , -- ADDR 388
			"00000000000000001000001101001111" , -- ADDR 389
			"00000000000000001011001111110001" , -- ADDR 390
			"00000000000000001100111100101110" , -- ADDR 391
			"00000000000000001000010110011101" , -- ADDR 392
			"00000000000000010010010110011110" , -- ADDR 393
			"00000000000000001101110100001010" , -- ADDR 394
			"00000000000000000111000010101100" , -- ADDR 395
			"00000000000000001101001101101000" , -- ADDR 396
			"00000000000000000110010110010000" , -- ADDR 397
			"00000000000000001100001001001011" , -- ADDR 398
			"00000000000000001101111110011101" , -- ADDR 399
			"00000000000000000100001011011101" , -- ADDR 400
			"00000000000000001100101111001101" , -- ADDR 401
			"00000000000000001100011110010000" , -- ADDR 402
			"00000000000000010100110001100000" , -- ADDR 403
			"00000000000000001101010110110100" , -- ADDR 404
			"00000000000000001110001011011110" , -- ADDR 405
			"00000000000000000111100101011000" , -- ADDR 406
			"00000000000000000110100100101110" , -- ADDR 407
			"00000000000000001111000110010111" , -- ADDR 408
			"00000000000000001010000000110100" , -- ADDR 409
			"00000000000000000011011111101110" , -- ADDR 410
			"00000000000000000010101011111000" , -- ADDR 411
			"00000000000000001001010010111111" , -- ADDR 412
			"00000000000000001101000111111111" , -- ADDR 413
			"00000000000000001001100110010111" , -- ADDR 414
			"00000000000000001101100111101001" , -- ADDR 415
			"00000000000000000101101100011100" , -- ADDR 416
			"00000000000000010011011000010011" , -- ADDR 417
			"00000000000000000100001011000000" , -- ADDR 418
			"00000000000000001101110111011110" , -- ADDR 419
			"00000000000000000101001110000010" , -- ADDR 420
			"00000000000000001110101010101011" , -- ADDR 421
			"00000000000000001001111000001100" , -- ADDR 422
			"00000000000000001101001011111001" , -- ADDR 423
			"00000000000000000010011100010000" , -- ADDR 424
			"00000000000000001111110000000010" , -- ADDR 425
			"00000000000000001101010111011001" , -- ADDR 426
			"00000000000000001101001001011100" , -- ADDR 427
			"00000000000000010000001110111011" , -- ADDR 428
			"00000000000000001110011011000100" , -- ADDR 429
			"00000000000000001011100100010101" , -- ADDR 430
			"00000000000000010010001100011101" , -- ADDR 431
			"00000000000000001111011001010111" , -- ADDR 432
			"00000000000000000110101010011111" , -- ADDR 433
			"00000000000000000100011010111111" , -- ADDR 434
			"00000000000000001001000010010110" , -- ADDR 435
			"00000000000000001000000101100001" , -- ADDR 436
			"00000000000000010001100110111101" , -- ADDR 437
			"00000000000000001111011001010111" , -- ADDR 438
			"00000000000000001101101010001010" , -- ADDR 439
			"00000000000000010100001110100111" , -- ADDR 440
			"00000000000000000110011111001011" , -- ADDR 441
			"00000000000000001110001010010000" , -- ADDR 442
			"00000000000000010001000101110000" , -- ADDR 443
			"00000000000000001101000000000110" , -- ADDR 444
			"00000000000000001001010110010000" , -- ADDR 445
			"00000000000000010010000100111001" , -- ADDR 446
			"00000000000000000111110010100010" , -- ADDR 447
			"00000000000000010010101000100010" , -- ADDR 448
			"00000000000000000110101001000011" , -- ADDR 449
			"00000000000000001110001110001001" , -- ADDR 450
			"00000000000000001010010000010000" , -- ADDR 451
			"00000000000000001110001100011010" , -- ADDR 452
			"00000000000000001111111001011011" , -- ADDR 453
			"00000000000000010010101111111000" , -- ADDR 454
			"00000000000000001000110011011000" , -- ADDR 455
			"00000000000000010111110110001001" , -- ADDR 456
			"00000000000000010011100010000000" , -- ADDR 457
			"00000000000000001000001111000110" , -- ADDR 458
			"00000000000000010011001110000001" , -- ADDR 459
			"00000000000000001000110110011001" , -- ADDR 460
			"00000000000000001100101101000110" , -- ADDR 461
			"00000000000000001110101010101011" , -- ADDR 462
			"00000000000000001100000011010110" , -- ADDR 463
			"00000000000000001111001011111001" , -- ADDR 464
			"00000000000000010110101110011110" , -- ADDR 465
			"00000000000000001110110000110001" , -- ADDR 466
			"00000000000000010010010011111111" , -- ADDR 467
			"00000000000000000100010001010101" , -- ADDR 468
			"00000000000000001010100001001001" , -- ADDR 469
			"00000000000000010010110110010001" , -- ADDR 470
			"00000000000000001010011111001001" , -- ADDR 471
			"00000000000000000110001110010111" , -- ADDR 472
			"00000000000000000101001110011001" , -- ADDR 473
			"00000000000000000101101100110001" , -- ADDR 474
			"00000000000000001101111110011101" , -- ADDR 475
			"00000000000000001101101100010000" , -- ADDR 476
			"00000000000000010001100101000111" , -- ADDR 477
			"00000000000000001001101010001000" , -- ADDR 478
			"00000000000000010001111101010001" , -- ADDR 479
			"00000000000000000001111101111110" , -- ADDR 480
			"00000000000000001100000111110001" , -- ADDR 481
			"00000000000000000001000101111000" , -- ADDR 482
			"00000000000000010010110011001110" , -- ADDR 483
			"00000000000000000110110010001001" , -- ADDR 484
			"00000000000000010001010110010111" , -- ADDR 485
			"00000000000000000011000011110010" , -- ADDR 486
			"00000000000000010001001000100010" , -- ADDR 487
			"00000000000000001110001100011010" , -- ADDR 488
			"00000000000000010001010010101111" , -- ADDR 489
			"00000000000000010100001110111001" , -- ADDR 490
			"00000000000000010001110011010110" , -- ADDR 491
			"00000000000000001111101001111101" , -- ADDR 492
			"00000000000000010001010101110100" , -- ADDR 493
			"00000000000000001110011010000000" , -- ADDR 494
			"00000000000000000111111110001010" , -- ADDR 495
			"00000000000000000110000100000111" , -- ADDR 496
			"00000000000000001001011001010100" , -- ADDR 497
			"00000000000000000110100110001011" , -- ADDR 498
			"00000000000000010000011000101111" , -- ADDR 499
			"00000000000000001101100000010101" , -- ADDR 500
			"00000000000000010001011000000001" , -- ADDR 501
			"00000000000000010101110011011100" , -- ADDR 502
			"00000000000000000011010100100001" , -- ADDR 503
			"00000000000000010001001000100010" , -- ADDR 504
			"00000000000000010011100001101101" , -- ADDR 505
			"00000000000000001111011000111000" , -- ADDR 506
			"00000000000000001100100011100110" , -- ADDR 507
			"00000000000000010011001110110100" , -- ADDR 508
			"00000000000000000101001111011111" , -- ADDR 509
			"00000000000000010100101111011111" , -- ADDR 510
			"00000000000000001010110001110011" , -- ADDR 511
			"00000000000000010001100101001110" , -- ADDR 512
			"00000000000000001110011010011010" , -- ADDR 513
			"00000000000000010000000110011011" , -- ADDR 514
			"00000000000000001111001011111001" , -- ADDR 515
			"00000000000000010011010100010000" , -- ADDR 516
			"00000000000000001100111100001000" , -- ADDR 517
			"00000000000000011010100000100001" , -- ADDR 518
			"00000000000000010101111011100100" , -- ADDR 519
			"00000000000000001100010001001001" , -- ADDR 520
			"00000000000000010100111100101010" , -- ADDR 521
			"00000000000000000111100101011000" , -- ADDR 522
			"00000000000000010000110111111100" , -- ADDR 523
			"00000000000000010010110101101010" , -- ADDR 524
			"00000000000000001011001000100111" , -- ADDR 525
			"00000000000000001110000110101111" , -- ADDR 526
			"00000000000000000110110101110010" , -- ADDR 527
			"00000000000000010100100001010110" , -- ADDR 528
			"00000000000000001001000100101010" , -- ADDR 529
			"00000000000000010001111010001011" , -- ADDR 530
			"00000000000000010001110111001100" , -- ADDR 531
			"00000000000000000011110100000100" , -- ADDR 532
			"00000000000000001010001010011101" , -- ADDR 533
			"00000000000000001111010111111000" , -- ADDR 534
			"00000000000000001001011110110001" , -- ADDR 535
			"00000000000000000100111010000100" , -- ADDR 536
			"00000000000000010000100101100101" , -- ADDR 537
			"00000000000000010010010000101001" , -- ADDR 538
			"00000000000000010001001001000110" , -- ADDR 539
			"00000000000000000110111010001110" , -- ADDR 540
			"00000000000000001101111110000011" , -- ADDR 541
			"00000000000000000011011010110000" , -- ADDR 542
			"00000000000000001011101110110100" , -- ADDR 543
			"00000000000000010100111011000111" , -- ADDR 544
			"00000000000000000111110100010000" , -- ADDR 545
			"00000000000000010100010100101001" , -- ADDR 546
			"00000000000000001010100100011010" , -- ADDR 547
			"00000000000000001000001011110110" , -- ADDR 548
			"00000000000000000100111100000000" , -- ADDR 549
			"00000000000000010110000110011001" , -- ADDR 550
			"00000000000000010100101000110000" , -- ADDR 551
			"00000000000000001111010010110010" , -- ADDR 552
			"00000000000000010001111011000010" , -- ADDR 553
			"00000000000000000101011101011001" , -- ADDR 554
			"00000000000000000010101110101100" , -- ADDR 555
			"00000000000000000110111010001110" , -- ADDR 556
			"00000000000000001000101010001100" , -- ADDR 557
			"00000000000000000100001100110101" , -- ADDR 558
			"00000000000000000101100000100001" , -- ADDR 559
			"00000000000000000101000001101111" , -- ADDR 560
			"00000000000000000100100011111010" , -- ADDR 561
			"00000000000000010000100110111101" , -- ADDR 562
			"00000000000000001100010110101110" , -- ADDR 563
			"00000000000000001111000010101100" , -- ADDR 564
			"00000000000000001101001101110001" , -- ADDR 565
			"00000000000000001100111111110011" , -- ADDR 566
			"00000000000000001010001001111001" , -- ADDR 567
			"00000000000000001011101001011011" , -- ADDR 568
			"00000000000000001001001101101000" , -- ADDR 569
			"00000000000000010001000011100001" , -- ADDR 570
			"00000000000000001100111010010111" , -- ADDR 571
			"00000000000000010001000000001010" , -- ADDR 572
			"00000000000000001111000011110101" , -- ADDR 573
			"00000000000000010001111101010001" , -- ADDR 574
			"00000000000000001001000010010110" , -- ADDR 575
			"00000000000000000011001011101110" , -- ADDR 576
			"00000000000000001000001000010110" , -- ADDR 577
			"00000000000000010000100100111001" , -- ADDR 578
			"00000000000000010011011111000100" , -- ADDR 579
			"00000000000000001110101111111111" , -- ADDR 580
			"00000000000000001111001100010001" , -- ADDR 581
			"00000000000000001100000001011100" , -- ADDR 582
			"00000000000000000100100000000111" , -- ADDR 583
			"00000000000000010100000110011001" , -- ADDR 584
			"00000000000000010101110001110010" , -- ADDR 585
			"00000000000000001000110100101011" , -- ADDR 586
			"00000000000000000101000010001000" , -- ADDR 587
			"00000000000000001010101100110101" , -- ADDR 588
			"00000000000000001111010111111000" , -- ADDR 589
			"00000000000000001101001010101111" , -- ADDR 590
			"00000000000000000110111010001110" , -- ADDR 591
			"00000000000000000111110100111110" , -- ADDR 592
			"00000000000000001001001001101011" , -- ADDR 593
			"00000000000000001110101000000100" , -- ADDR 594
			"00000000000000010000110101100100" , -- ADDR 595
			"00000000000000000110110010001001" , -- ADDR 596
			"00000000000000001000011011011101" , -- ADDR 597
			"00000000000000000111111110001010" , -- ADDR 598
			"00000000000000001100110110010111" , -- ADDR 599
			"00000000000000010000110111111100" , -- ADDR 600
			"00000000000000010000001111100000" , -- ADDR 601
			"00000000000000001110011101011100" , -- ADDR 602
			"00000000000000001111101101011111" , -- ADDR 603
			"00000000000000001010111111001000" , -- ADDR 604
			"00000000000000001111111100011011" , -- ADDR 605
			"00000000000000001011000001111001" , -- ADDR 606
			"00000000000000001100001010011100" , -- ADDR 607
			"00000000000000000110000111100100" , -- ADDR 608
			"00000000000000000110111010001110" , -- ADDR 609
			"00000000000000001101101111101111" , -- ADDR 610
			"00000000000000001001111010100000" , -- ADDR 611
			"00000000000000000100001011000000" , -- ADDR 612
			"00000000000000001000110000000111" , -- ADDR 613
			"00000000000000001110010111000110" , -- ADDR 614
			"00000000000000001101000111010000" , -- ADDR 615
			"00000000000000000111101010011001" , -- ADDR 616
			"00000000000000001001001001000011" , -- ADDR 617
			"00000000000000001000010100001011" , -- ADDR 618
			"00000000000000001100001101011010" , -- ADDR 619
			"00000000000000001111000101001110" , -- ADDR 620
			"00000000000000001111101100100000" , -- ADDR 621
			"00000000000000000101111000010011" , -- ADDR 622
			"00000000000000001001000010001000" , -- ADDR 623
			"00000000000000010010011000010110" , -- ADDR 624
			"00000000000000000010001101011111" , -- ADDR 625
			"00000000000000000100101100100011" , -- ADDR 626
			"00000000000000000001011011000111" , -- ADDR 627
			"00000000000000000011100011100000" , -- ADDR 628
			"00000000000000001000010110000000" , -- ADDR 629
			"00000000000000010100000010011001" , -- ADDR 630
			"00000000000000000110100100101110" , -- ADDR 631
			"00000000000000001011100110011110" , -- ADDR 632
			"00000000000000000011111100011011" , -- ADDR 633
			"00000000000000001001110001011001" , -- ADDR 634
			"00000000000000000011100110101101" , -- ADDR 635
			"00000000000000001100100100010110" , -- ADDR 636
			"00000000000000001010100000100110" , -- ADDR 637
			"00000000000000001001000100000001" , -- ADDR 638
			"00000000000000001011011001001101" , -- ADDR 639
			"00000000000000000111000111100011" , -- ADDR 640
			"00000000000000000111110100000000" , -- ADDR 641
			"00000000000000000111110100010000" , -- ADDR 642
			"00000000000000001011110011110110" , -- ADDR 643
			"00000000000000001011000010000100" , -- ADDR 644
			"00000000000000001100001100001010" , -- ADDR 645
			"00000000000000001000001000010110" , -- ADDR 646
			"00000000000000010001110001001100" , -- ADDR 647
			"00000000000000010101101010011010" , -- ADDR 648
			"00000000000000010101111110101100" , -- ADDR 649
			"00000000000000001100101111101010" , -- ADDR 650
			"00000000000000001100110110010111" , -- ADDR 651
			"00000000000000010001010010101111" , -- ADDR 652
			"00000000000000010111001001011010" , -- ADDR 653
			"00000000000000010110101101001101" , -- ADDR 654
			"00000000000000001001100011001011" , -- ADDR 655
			"00000000000000010000110111001001" , -- ADDR 656
			"00000000000000001110111100000100" , -- ADDR 657
			"00000000000000010101101011000001" , -- ADDR 658
			"00000000000000010000100110100111" , -- ADDR 659
			"00000000000000011000000111111101" , -- ADDR 660
			"00000000000000010001010010110110" , -- ADDR 661
			"00000000000000010110111111011111" , -- ADDR 662
			"00000000000000010001111000011110" , -- ADDR 663
			"00000000000000010101010101000111" , -- ADDR 664
			"00000000000000010010100010110010" , -- ADDR 665
			"00000000000000010011111011001001" , -- ADDR 666
			"00000000000000000110000001111010" , -- ADDR 667
			"00000000000000001001011010111100" , -- ADDR 668
			"00000000000000010101100111110110" , -- ADDR 669
			"00000000000000001111101100000001" , -- ADDR 670
			"00000000000000001010001001111001" , -- ADDR 671
			"00000000000000010000101001011000" , -- ADDR 672
			"00000000000000001101111010110001" , -- ADDR 673
			"00000000000000001110100000101111" , -- ADDR 674
			"00000000000000001110110000011000" , -- ADDR 675
			"00000000000000010000110011010011" , -- ADDR 676
			"00000000000000001101110110010111" , -- ADDR 677
			"00000000000000010001111011000010" , -- ADDR 678
			"00000000000000001111011011011110" , -- ADDR 679
			"00000000000000010001111000011110" , -- ADDR 680
			"00000000000000001100101001001100" , -- ADDR 681
			"00000000000000000010010000000100" , -- ADDR 682
			"00000000000000011010000010101100" , -- ADDR 683
			"00000000000000001000010011010000" , -- ADDR 684
			"00000000000000000100011001010000" , -- ADDR 685
			"00000000000000000111111000110111" , -- ADDR 686
			"00000000000000001100011000000111" , -- ADDR 687
			"00000000000000000101001011011101" , -- ADDR 688
			"00000000000000011011111000011010" , -- ADDR 689
			"00000000000000000010010000000100" , -- ADDR 690
			"00000000000000010100011001011010" , -- ADDR 691
			"00000000000000001010000111011101" , -- ADDR 692
			"00000000000000010010000100010000" , -- ADDR 693
			"00000000000000000110101001000011" , -- ADDR 694
			"00000000000000001101011010000110" , -- ADDR 695
			"00000000000000000111100101011000" , -- ADDR 696
			"00000000000000010001101000111010" , -- ADDR 697
			"00000000000000000101111000010011" , -- ADDR 698
			"00000000000000000010110110001110" , -- ADDR 699
			"00000000000000010000100000010010" , -- ADDR 700
			"00000000000000000010000101100000" , -- ADDR 701
			"00000000000000010001001001000110" , -- ADDR 702
			"00000000000000010010101101101111" , -- ADDR 703
			"00000000000000010011010011100100" , -- ADDR 704
			"00000000000000001111100110010011" , -- ADDR 705
			"00000000000000001101100010010100" , -- ADDR 706
			"00000000000000010000001011100000" , -- ADDR 707
			"00000000000000001011111010111010" , -- ADDR 708
			"00000000000000000100101111011000" , -- ADDR 709
			"00000000000000001001111001001010" , -- ADDR 710
			"00000000000000001111111011100101" , -- ADDR 711
			"00000000000000001110101000000100" , -- ADDR 712
			"00000000000000000001111101111110" , -- ADDR 713
			"00000000000000001100101010110110" , -- ADDR 714
			"00000000000000001100111100101110" , -- ADDR 715
			"00000000000000001111101001000110" , -- ADDR 716
			"00000000000000001011111001111101" , -- ADDR 717
			"00000000000000010000010010101011" , -- ADDR 718
			"00000000000000001010010000011100" , -- ADDR 719
			"00000000000000001110111100100101" , -- ADDR 720
			"00000000000000001111111010101000" , -- ADDR 721
			"00000000000000001101010100111101" , -- ADDR 722
			"00000000000000001111110001111101" , -- ADDR 723
			"00000000000000001100000111110001" , -- ADDR 724
			"00000000000000000010011001111001" , -- ADDR 725
			"00000000000000000010000000110110" , -- ADDR 726
			"00000000000000010010001111010010" , -- ADDR 727
			"00000000000000001110111100100101" , -- ADDR 728
			"00000000000000001001000101100000" , -- ADDR 729
			"00000000000000001101011010000110" , -- ADDR 730
			"00000000000000001001010110000011" , -- ADDR 731
			"00000000000000001000010110011101" , -- ADDR 732
			"00000000000000000110111000010010" , -- ADDR 733
			"00000000000000001001000100101010" , -- ADDR 734
			"00000000000000000101101110000111" , -- ADDR 735
			"00000000000000001001110100100000" , -- ADDR 736
			"00000000000000001010001010011101" , -- ADDR 737
			"00000000000000001011010001011110" , -- ADDR 738
			"00000000000000001010111010010000" , -- ADDR 739
			"00000000000000000111000010101100" , -- ADDR 740
			"00000000000000010010000101001101" , -- ADDR 741
			"00000000000000000110110001010011" , -- ADDR 742
			"00000000000000000110001011100110" , -- ADDR 743
			"00000000000000000011101110100000" , -- ADDR 744
			"00000000000000000111001101101011" , -- ADDR 745
			"00000000000000000100101111011000" , -- ADDR 746
			"00000000000000010011111110101011" , -- ADDR 747
			"00000000000000000110011100110100" , -- ADDR 748
			"00000000000000001110110011111111" , -- ADDR 749
			"00000000000000001000111000000111" , -- ADDR 750
			"00000000000000001110000101100001" , -- ADDR 751
			"00000000000000000010001100101000" , -- ADDR 752
			"00000000000000000111101010011001" , -- ADDR 753
			"00000000000000000110000010100011" , -- ADDR 754
			"00000000000000001101000011110000" , -- ADDR 755
			"00000000000000001100111010111100" , -- ADDR 756
			"00000000000000001000000111011010" , -- ADDR 757
			"00000000000000001011101010010000" , -- ADDR 758
			"00000000000000000110001110010111" , -- ADDR 759
			"00000000000000001001000101100000" , -- ADDR 760
			"00000000000000001111101101011111" , -- ADDR 761
			"00000000000000010001000010110110" , -- ADDR 762
			"00000000000000010100110010100111" , -- ADDR 763
			"00000000000000001001011111111110" , -- ADDR 764
			"00000000000000000101001000100000" , -- ADDR 765
			"00000000000000010000101110011001" , -- ADDR 766
			"00000000000000001100111011011001" , -- ADDR 767
			"00000000000000001110100100010010" , -- ADDR 768
			"00000000000000010110100011101100" , -- ADDR 769
			"00000000000000010001000101110111" , -- ADDR 770
			"00000000000000000100101010100001" , -- ADDR 771
			"00000000000000000010110110111001" , -- ADDR 772
			"00000000000000001001111110010101" , -- ADDR 773
			"00000000000000011011000000101011" , -- ADDR 774
			"00000000000000010010001100110001" , -- ADDR 775
			"00000000000000010111011010001000" , -- ADDR 776
			"00000000000000010011010010011110" , -- ADDR 777
			"00000000000000000000011111010000" , -- ADDR 778
			"00000000000000010110011100010100" , -- ADDR 779
			"00000000000000000001011000011001" , -- ADDR 780
			"00000000000000001111101011000011" , -- ADDR 781
			"00000000000000010000110010111101" , -- ADDR 782
			"00000000000000010001010001000101" , -- ADDR 783
			"00000000000000000100011001101100" , -- ADDR 784
			"00000000000000000011001011101110" , -- ADDR 785
			"00000000000000000111101001011001" , -- ADDR 786
			"00000000000000000010110010001010" , -- ADDR 787
			"00000000000000011000101100010011" , -- ADDR 788
			"00000000000000010110111101000101" , -- ADDR 789
			"00000000000000001110011011010101" , -- ADDR 790
			"00000000000000001110001001110110" , -- ADDR 791
			"00000000000000010000101000000000" , -- ADDR 792
			"00000000000000010011001001100011" , -- ADDR 793
			"00000000000000011001001000011110" , -- ADDR 794
			"00000000000000011000110111110000" , -- ADDR 795
			"00000000000000000101001011000110" , -- ADDR 796
			"00000000000000010010110101101010" , -- ADDR 797
			"00000000000000010100011110010111" , -- ADDR 798
			"00000000000000001001110101110111" , -- ADDR 799
			"00000000000000001101100001000010" , -- ADDR 800
			"00000000000000001100000111110001" , -- ADDR 801
			"00000000000000001000111000110001" , -- ADDR 802
			"00000000000000010010111001100110" , -- ADDR 803
			"00000000000000010101010100011001" , -- ADDR 804
			"00000000000000001111110000110000" , -- ADDR 805
			"00000000000000001000010000101110" , -- ADDR 806
			"00000000000000000111101110000111" , -- ADDR 807
			"00000000000000000011111110010111" , -- ADDR 808
			"00000000000000001110010010011011" , -- ADDR 809
			"00000000000000010110101010110001" , -- ADDR 810
			"00000000000000010101001100100110" , -- ADDR 811
			"00000000000000000101011000000111" , -- ADDR 812
			"00000000000000010000111101010110" , -- ADDR 813
			"00000000000000001111000101110110" , -- ADDR 814
			"00000000000000000110001011100110" , -- ADDR 815
			"00000000000000010001100110101111" , -- ADDR 816
			"00000000000000010011010001001100" , -- ADDR 817
			"00000000000000000001111010000010" , -- ADDR 818
			"00000000000000000001100010110101" , -- ADDR 819
			"00000000000000001110001001111111" , -- ADDR 820
			"00000000000000010100010101011111" , -- ADDR 821
			"00000000000000001000110100011101" , -- ADDR 822
			"00000000000000000111110111111001" , -- ADDR 823
			"00000000000000001001010101000010" , -- ADDR 824
			"00000000000000000001110001110000" , -- ADDR 825
			"00000000000000001100010000100010" , -- ADDR 826
			"00000000000000010000001000110010" , -- ADDR 827
			"00000000000000010011100010111000" , -- ADDR 828
			"00000000000000001101010001101010" , -- ADDR 829
			"00000000000000001110001010010000" , -- ADDR 830
			"00000000000000000110000111111000" , -- ADDR 831
			"00000000000000001000010011011111" , -- ADDR 832
			"00000000000000000011011001101000" , -- ADDR 833
			"00000000000000010101010001011100" , -- ADDR 834
			"00000000000000000010100000111000" , -- ADDR 835
			"00000000000000010100000001010000" , -- ADDR 836
			"00000000000000000101010110101100" , -- ADDR 837
			"00000000000000001111101101111110" , -- ADDR 838
			"00000000000000001100011011110011" , -- ADDR 839
			"00000000000000010100011111011110" , -- ADDR 840
			"00000000000000010110001110101001" , -- ADDR 841
			"00000000000000010010101110010000" , -- ADDR 842
			"00000000000000010010000001100000" , -- ADDR 843
			"00000000000000001101111011101110" , -- ADDR 844
			"00000000000000001011000001000010" , -- ADDR 845
			"00000000000000000111101110000111" , -- ADDR 846
			"00000000000000000110110101110010" , -- ADDR 847
			"00000000000000000111110100010000" , -- ADDR 848
			"00000000000000000011110100000100" , -- ADDR 849
			"00000000000000001100110000010000" , -- ADDR 850
			"00000000000000001001100011001011" , -- ADDR 851
			"00000000000000010010110110110001" , -- ADDR 852
			"00000000000000010100010111101111" , -- ADDR 853
			"00000000000000000110010110100011" , -- ADDR 854
			"00000000000000010001100001101000" , -- ADDR 855
			"00000000000000010011001000110110" , -- ADDR 856
			"00000000000000001111001011011001" , -- ADDR 857
			"00000000000000001101100100011011" , -- ADDR 858
			"00000000000000010001011110100101" , -- ADDR 859
			"00000000000000001000010011011111" , -- ADDR 860
			"00000000000000010011111011001001" , -- ADDR 861
			"00000000000000001110000101100001" , -- ADDR 862
			"00000000000000010010011110111110" , -- ADDR 863
			"00000000000000010001000111001101" , -- ADDR 864
			"00000000000000001111010011011010" , -- ADDR 865
			"00000000000000001011111110010001" , -- ADDR 866
			"00000000000000010001000000001010" , -- ADDR 867
			"00000000000000001111100100101101" , -- ADDR 868
			"00000000000000011010001010110011" , -- ADDR 869
			"00000000000000010101011001110000" , -- ADDR 870
			"00000000000000001110100111000001" , -- ADDR 871
			"00000000000000010011101101010010" , -- ADDR 872
			"00000000000000000100101111011000" , -- ADDR 873
			"00000000000000010011100110011001" , -- ADDR 874
			"00000000000000010101100011100111" , -- ADDR 875
			"00000000000000001100011100101110" , -- ADDR 876
			"00000000000000001110011101100101" , -- ADDR 877
			"00000000000000000111110010100010" , -- ADDR 878
			"00000000000000000101101010011011" , -- ADDR 879
			"00000000000000001111110111101000" , -- ADDR 880
			"00000000000000010000101101011111" , -- ADDR 881
			"00000000000000000110000100000111" , -- ADDR 882
			"00000000000000001010001100101101" , -- ADDR 883
			"00000000000000000000111000010110" , -- ADDR 884
			"00000000000000011000110011011101" , -- ADDR 885
			"00000000000000001001101110000100" , -- ADDR 886
			"00000000000000010011101110100010" , -- ADDR 887
			"00000000000000001011100110110011" , -- ADDR 888
			"00000000000000001001111100001111" , -- ADDR 889
			"00000000000000010000011010000001" , -- ADDR 890
			"00000000000000001000001101001111" , -- ADDR 891
			"00000000000000001000111000110001" , -- ADDR 892
			"00000000000000010010010100010011" , -- ADDR 893
			"00000000000000010000111100110010" , -- ADDR 894
			"00000000000000000111000101001000" , -- ADDR 895
			"00000000000000001100010100101110" , -- ADDR 896
			"00000000000000001101000111010000" , -- ADDR 897
			"00000000000000000111101000001001" , -- ADDR 898
			"00000000000000010111001011011001" , -- ADDR 899
			"00000000000000010100101000110110" , -- ADDR 900
			"00000000000000001011000010000100" , -- ADDR 901
			"00000000000000001001010110000011" , -- ADDR 902
			"00000000000000001101110000101101" , -- ADDR 903
			"00000000000000001110001011000100" , -- ADDR 904
			"00000000000000010110111011110101" , -- ADDR 905
			"00000000000000010101010010100001" , -- ADDR 906
			"00000000000000001011010101000000" , -- ADDR 907
			"00000000000000010110000110111010" , -- ADDR 908
			"00000000000000001011110010000100" , -- ADDR 909
			"00000000000000001101111110011101" , -- ADDR 910
			"00000000000000010001101101010101" , -- ADDR 911
			"00000000000000001110010000110101" , -- ADDR 912
			"00000000000000001001101000100011" , -- ADDR 913
			"00000000000000010100110000100000" , -- ADDR 914
			"00000000000000001100001110101010" , -- ADDR 915
			"00000000000000010011101110101000" , -- ADDR 916
			"00000000000000000001101000110100" , -- ADDR 917
			"00000000000000001100111111110011" , -- ADDR 918
			"00000000000000000101110000110001" , -- ADDR 919
			"00000000000000010000001000010100" , -- ADDR 920
			"00000000000000010100110111110101" , -- ADDR 921
			"00000000000000010110001010101100" , -- ADDR 922
			"00000000000000000101000010001000" , -- ADDR 923
			"00000000000000010111011110010111" , -- ADDR 924
			"00000000000000010011111111110100" , -- ADDR 925
			"00000000000000000101101011011011" , -- ADDR 926
			"00000000000000010100111011001101" , -- ADDR 927
			"00000000000000001110110000011000" , -- ADDR 928
			"00000000000000000111101010011001" , -- ADDR 929
			"00000000000000001001011011001001" , -- ADDR 930
			"00000000000000001110010010011011" , -- ADDR 931
			"00000000000000001100101111001101" , -- ADDR 932
			"00000000000000010000010101001000" , -- ADDR 933
			"00000000000000010110000000011011" , -- ADDR 934
			"00000000000000001101101100010000" , -- ADDR 935
			"00000000000000000110011000111101" , -- ADDR 936
			"00000000000000000010100011001000" , -- ADDR 937
			"00000000000000001100100110101000" , -- ADDR 938
			"00000000000000010111110010001001" , -- ADDR 939
			"00000000000000010011010001001100" , -- ADDR 940
			"00000000000000010101000100111011" , -- ADDR 941
			"00000000000000010011101010001011" , -- ADDR 942
			"00000000000000000101001011011101" , -- ADDR 943
			"00000000000000010101011111010111" , -- ADDR 944
			"00000000000000000110001001011011" , -- ADDR 945
			"00000000000000001111110111101000" , -- ADDR 946
			"00000000000000001100100110101000" , -- ADDR 947
			"00000000000000001101110100011100" , -- ADDR 948
			"00000000000000001001010110111000" , -- ADDR 949
			"00000000000000000011001000000110" , -- ADDR 950
			"00000000000000000010111100001010" , -- ADDR 951
			"00000000000000000101000001101111" , -- ADDR 952
			"00000000000000010101010000110100" , -- ADDR 953
			"00000000000000010011111110110001" , -- ADDR 954
			"00000000000000001100111101011101" , -- ADDR 955
			"00000000000000001101100000011110" , -- ADDR 956
			"00000000000000001110100000101111" , -- ADDR 957
			"00000000000000010001110111010011" , -- ADDR 958
			"00000000000000010101111111000010" , -- ADDR 959
			"00000000000000010110011001110001" , -- ADDR 960
			"00000000000000000001011111000011" , -- ADDR 961
			"00000000000000001101111110110111" , -- ADDR 962
			"00000000000000010101100101000111" , -- ADDR 963
			"00000000000000000101010110101100" , -- ADDR 964
			"00000000000000001000101000001101" , -- ADDR 965
			"00000000000000001000001101000001" , -- ADDR 966
			"00000000000000000110110101110010" , -- ADDR 967
			"00000000000000001110011101000011" , -- ADDR 968
			"00000000000000010110110100100000" , -- ADDR 969
			"00000000000000001010110101100001" , -- ADDR 970
			"00000000000000001010111000001001" , -- ADDR 971
			"00000000000000000011000110111000" , -- ADDR 972
			"00000000000000000110111010001110" , -- ADDR 973
			"00000000000000001010001100101101" , -- ADDR 974
			"00000000000000010011011110001100" , -- ADDR 975
			"00000000000000010000111100110010" , -- ADDR 976
			"00000000000000000111011011001110" , -- ADDR 977
			"00000000000000001011111011000100" , -- ADDR 978
			"00000000000000001010000000101000" , -- ADDR 979
			"00000000000000000111001011100011" , -- ADDR 980
			"00000000000000001100110001100110" , -- ADDR 981
			"00000000000000010001101101110000" , -- ADDR 982
			"00000000000000000110011101101100" , -- ADDR 983
			"00000000000000000110101000011110" , -- ADDR 984
			"00000000000000000110111100011011" , -- ADDR 985
			"00000000000000001100101100101010" , -- ADDR 986
			"00000000000000001001111000110001" , -- ADDR 987
			"00000000000000000011100001010110" , -- ADDR 988
			"00000000000000001100110001111001" , -- ADDR 989
			"00000000000000001110100001011001" , -- ADDR 990
			"00000000000000001101101111101111" , -- ADDR 991
			"00000000000000001010100110011001" , -- ADDR 992
			"00000000000000001100001100111100" , -- ADDR 993
			"00000000000000000110110011010001" , -- ADDR 994
			"00000000000000001010100000100110" , -- ADDR 995
			"00000000000000010001001000100010" , -- ADDR 996
			"00000000000000001000101000001101" , -- ADDR 997
			"00000000000000010000100000101000" , -- ADDR 998
			"00000000000000001000001111000110" , -- ADDR 999
			"00000000000000000110111001111100" , -- ADDR 1000
			"00000000000000000011101110100000" , -- ADDR 1001
			"00000000000000010010010011111111" , -- ADDR 1002
			"00000000000000010000111101010110" , -- ADDR 1003
			"00000000000000001011111000010110" , -- ADDR 1004
			"00000000000000001110000111001001" , -- ADDR 1005
			"00000000000000001000101111000001" , -- ADDR 1006
			"00000000000000000110011010001001" , -- ADDR 1007
			"00000000000000000011011111101110" , -- ADDR 1008
			"00000000000000000101100111101110" , -- ADDR 1009
			"00000000000000000001000101111000" , -- ADDR 1010
			"00000000000000000101000101001001" , -- ADDR 1011
			"00000000000000001000101100011001" , -- ADDR 1012
			"00000000000000001000001100000101" , -- ADDR 1013
			"00000000000000001100111110010101" , -- ADDR 1014
			"00000000000000001011100101000000" , -- ADDR 1015
			"00000000000000001101110000100100" , -- ADDR 1016
			"00000000000000001010000000110100" , -- ADDR 1017
			"00000000000000001010101010001010" , -- ADDR 1018
			"00000000000000000111000111100011" , -- ADDR 1019
			"00000000000000000111110111111001" , -- ADDR 1020
			"00000000000000001000110011011000" , -- ADDR 1021
			"00000000000000001111101110010101" , -- ADDR 1022
			"00000000000000001011001011100001" , -- ADDR 1023
			"00000000000000001101011011100001" , -- ADDR 1024
			"00000000000000001011101000111100" , -- ADDR 1025
			"00000000000000001110001001111111" , -- ADDR 1026
			"00000000000000000110101010110001" , -- ADDR 1027
			"00000000000000000110011100110100" , -- ADDR 1028
			"00000000000000001000111000110001" , -- ADDR 1029
			"00000000000000001100110010110010" , -- ADDR 1030
			"00000000000000010001100101001110" , -- ADDR 1031
			"00000000000000001100110001100110" , -- ADDR 1032
			"00000000000000001011011001100010" , -- ADDR 1033
			"00000000000000001010111000110110" , -- ADDR 1034
			"00000000000000000100010111100001" , -- ADDR 1035
			"00000000000000010000010010010100" , -- ADDR 1036
			"00000000000000010001111110000000" , -- ADDR 1037
			"00000000000000000110000010100011" , -- ADDR 1038
			"00000000000000001001101000100011" , -- ADDR 1039
			"00000000000000001001110010110000" , -- ADDR 1040
			"00000000000000001000010010100100" , -- ADDR 1041
			"00000000000000001011101110001010" , -- ADDR 1042
			"00000000000000000110111111101101" , -- ADDR 1043
			"00000000000000010001000010001011" , -- ADDR 1044
			"00000000000000000111000110001101" , -- ADDR 1045
			"00000000000000001011111110010001" , -- ADDR 1046
			"00000000000000000110111100101100" , -- ADDR 1047
			"00000000000000001101011010000110" , -- ADDR 1048
			"00000000000000001001100100110001" , -- ADDR 1049
			"00000000000000001100001101010000" , -- ADDR 1050
			"00000000000000000011001011001000" , -- ADDR 1051
			"00000000000000001100010001110001" , -- ADDR 1052
			"00000000000000001010000010010110" , -- ADDR 1053
			"00000000000000001101000001011011" , -- ADDR 1054
			"00000000000000001110011010000000" , -- ADDR 1055
			"00000000000000001011100101000000" , -- ADDR 1056
			"00000000000000001010001001111001" , -- ADDR 1057
			"00000000000000001111100001010001" , -- ADDR 1058
			"00000000000000001100111001000010" , -- ADDR 1059
			"00000000000000000011011100111110" , -- ADDR 1060
			"00000000000000000001100100000011" , -- ADDR 1061
			"00000000000000000110000110101000" , -- ADDR 1062
			"00000000000000000110101001000011" , -- ADDR 1063
			"00000000000000001111001011011001" , -- ADDR 1064
			"00000000000000001101100010010100" , -- ADDR 1065
			"00000000000000001011010000010010" , -- ADDR 1066
			"00000000000000010000101110111110" , -- ADDR 1067
			"00000000000000001001010001111101" , -- ADDR 1068
			"00000000000000001010111111001000" , -- ADDR 1069
			"00000000000000001101101100010000" , -- ADDR 1070
			"00000000000000001001100100100101" , -- ADDR 1071
			"00000000000000000110010101010110" , -- ADDR 1072
			"00000000000000001110101000000100" , -- ADDR 1073
			"00000000000000001010111000110110" , -- ADDR 1074
			"00000000000000001111001010110001" , -- ADDR 1075
			"00000000000000000111000101001000" , -- ADDR 1076
			"00000000000000001011010110110111" , -- ADDR 1077
			"00000000000000001001010110000011" , -- ADDR 1078
			"00000000000000001010101100110101" , -- ADDR 1079
			"00000000000000001101001101000011" , -- ADDR 1080
			"00000000000000001111011011011110" , -- ADDR 1081
			"00000000000000000111110011010001" , -- ADDR 1082
			"00000000000000010100100010110101" , -- ADDR 1083
			"00000000000000010000001000010100" , -- ADDR 1084
			"00000000000000000110110000001011" , -- ADDR 1085
			"00000000000000001111101110010101" , -- ADDR 1086
			"00000000000000000111000101001000" , -- ADDR 1087
			"00000000000000001011110100000000" , -- ADDR 1088
			"00000000000000001101110000000001" , -- ADDR 1089
			"00000000000000001010111000110110" , -- ADDR 1090
			"00000000000000001111110001110110" , -- ADDR 1091
			"00000000000000001010010010101010" , -- ADDR 1092
			"00000000000000001110100001110010" , -- ADDR 1093
			"00000000000000000100111000111001" , -- ADDR 1094
			"00000000000000010101111011110100" , -- ADDR 1095
			"00000000000000000100000101111011" , -- ADDR 1096
			"00000000000000010000010100100011" , -- ADDR 1097
			"00000000000000000110010011001111" , -- ADDR 1098
			"00000000000000001111000010101100" , -- ADDR 1099
			"00000000000000001011110010001110" , -- ADDR 1100
			"00000000000000001101011010000110" , -- ADDR 1101
			"00000000000000000100110111010101" , -- ADDR 1102
			"00000000000000010010010011111000" , -- ADDR 1103
			"00000000000000010000000001010100" , -- ADDR 1104
			"00000000000000001100101101110110" , -- ADDR 1105
			"00000000000000010001000000001010" , -- ADDR 1106
			"00000000000000010000000101000000" , -- ADDR 1107
			"00000000000000001100001100111100" , -- ADDR 1108
			"00000000000000010100110101010001" , -- ADDR 1109
			"00000000000000010010000000011100" , -- ADDR 1110
			"00000000000000001001010101000010" , -- ADDR 1111
			"00000000000000000111000110001101" , -- ADDR 1112
			"00000000000000001011101110001010" , -- ADDR 1113
			"00000000000000001010100001001001" , -- ADDR 1114
			"00000000000000010100001100010110" , -- ADDR 1115
			"00000000000000010001110100101111" , -- ADDR 1116
			"00000000000000001110111101101110" , -- ADDR 1117
			"00000000000000010110101101111000" , -- ADDR 1118
			"00000000000000000110000111111000" , -- ADDR 1119
			"00000000000000010000001000010100" , -- ADDR 1120
			"00000000000000010011010011100100" , -- ADDR 1121
			"00000000000000001111010010111010" , -- ADDR 1122
			"00000000000000001011010010010100" , -- ADDR 1123
			"00000000000000010100101010100110" , -- ADDR 1124
			"00000000000000000110110000001011" , -- ADDR 1125
			"00000000000000010100111101111100" , -- ADDR 1126
			"00000000000000000110011000111101" , -- ADDR 1127
			"00000000000000001111111001011011" , -- ADDR 1128
			"00000000000000001010100110011001" , -- ADDR 1129
			"00000000000000010000101000111010" , -- ADDR 1130
			"00000000000000010010100010110010" , -- ADDR 1131
			"00000000000000010101011010001101" , -- ADDR 1132
			"00000000000000001001010110000011" , -- ADDR 1133
			"00000000000000011001111000111010" , -- ADDR 1134
			"00000000000000010101101111010101" , -- ADDR 1135
			"00000000000000001001001011010110" , -- ADDR 1136
			"00000000000000010101101011000001" , -- ADDR 1137
			"00000000000000001011010110010111" , -- ADDR 1138
			"00000000000000001100111000100101" , -- ADDR 1139
			"00000000000000001110110001110011" , -- ADDR 1140
			"00000000000000001101001100010101" , -- ADDR 1141
			"00000000000000010001111010000100" , -- ADDR 1142
			"00000000000000010101010001101000" , -- ADDR 1143
			"00000000000000001110111111011000" , -- ADDR 1144
			"00000000000000001101110001110100" , -- ADDR 1145
			"00000000000000000111011000011000" , -- ADDR 1146
			"00000000000000001000000011011001" , -- ADDR 1147
			"00000000000000000100101100001001" , -- ADDR 1148
			"00000000000000010111000010011110" , -- ADDR 1149
			"00000000000000000001110001110000" , -- ADDR 1150
			"00000000000000010101110010110101" , -- ADDR 1151
			"00000000000000000111000111100011" , -- ADDR 1152
			"00000000000000010000101100111011" , -- ADDR 1153
			"00000000000000001101010110010000" , -- ADDR 1154
			"00000000000000010110010000101101" , -- ADDR 1155
			"00000000000000010111111101001111" , -- ADDR 1156
			"00000000000000010100010011110011" , -- ADDR 1157
			"00000000000000010011110010011001" , -- ADDR 1158
			"00000000000000001101111001011001" , -- ADDR 1159
			"00000000000000001011000011111110" , -- ADDR 1160
			"00000000000000001001001111011111" , -- ADDR 1161
			"00000000000000001000100011000110" , -- ADDR 1162
			"00000000000000001000111101101011" , -- ADDR 1163
			"00000000000000000100110100001011" , -- ADDR 1164
			"00000000000000001100100011011100" , -- ADDR 1165
			"00000000000000001001000101100000" , -- ADDR 1166
			"00000000000000010100100001111111" , -- ADDR 1167
			"00000000000000010101010010100111" , -- ADDR 1168
			"00000000000000000111000111000000" , -- ADDR 1169
			"00000000000000010011000000111101" , -- ADDR 1170
			"00000000000000010100011010101110" , -- ADDR 1171
			"00000000000000010000100011000011" , -- ADDR 1172
			"00000000000000001111001101010010" , -- ADDR 1173
			"00000000000000010010010011010111" , -- ADDR 1174
			"00000000000000001000111010010001" , -- ADDR 1175
			"00000000000000010101000100001100" , -- ADDR 1176
			"00000000000000001111110101110101" , -- ADDR 1177
			"00000000000000010100000100011001" , -- ADDR 1178
			"00000000000000010010111000111001" , -- ADDR 1179
			"00000000000000010000100000010010" , -- ADDR 1180
			"00000000000000001100000111111011" , -- ADDR 1181
			"00000000000000010001100101000111" , -- ADDR 1182
			"00000000000000010001010110010111" , -- ADDR 1183
			"00000000000000011011011010100110" , -- ADDR 1184
			"00000000000000010110100111110101" , -- ADDR 1185
			"00000000000000010000011000001010" , -- ADDR 1186
			"00000000000000010100101101001100" , -- ADDR 1187
			"00000000000000000101100100010100" , -- ADDR 1188
			"00000000000000010101011000000100" , -- ADDR 1189
			"00000000000000010111010101001111" , -- ADDR 1190
			"00000000000000001101110100011100" , -- ADDR 1191
			"00000000000000001110100010011100" , -- ADDR 1192
			"00000000000000010000000110000100" , -- ADDR 1193
			"00000000000000001010000101111100" , -- ADDR 1194
			"00000000000000001111101001001110" , -- ADDR 1195
			"00000000000000001000010100001011" , -- ADDR 1196
			"00000000000000001110000001101110" , -- ADDR 1197
			"00000000000000010001011011111101" , -- ADDR 1198
			"00000000000000001011110010000100" , -- ADDR 1199
			"00000000000000010001001010010100" , -- ADDR 1200
			"00000000000000001011100101001010" , -- ADDR 1201
			"00000000000000000011100001010110" , -- ADDR 1202
			"00000000000000000000001111101000" , -- ADDR 1203
			"00000000000000010011011011111100" , -- ADDR 1204
			"00000000000000010000101010010010" , -- ADDR 1205
			"00000000000000001010111010110001" , -- ADDR 1206
			"00000000000000001110110000011000" , -- ADDR 1207
			"00000000000000000111101000001001" , -- ADDR 1208
			"00000000000000000110011010001001" , -- ADDR 1209
			"00000000000000000110011101101100" , -- ADDR 1210
			"00000000000000001000101101101101" , -- ADDR 1211
			"00000000000000000100100110110100" , -- ADDR 1212
			"00000000000000001000011101011111" , -- ADDR 1213
			"00000000000000001000010011010000" , -- ADDR 1214
			"00000000000000001001010011100110" , -- ADDR 1215
			"00000000000000001100100110011110" , -- ADDR 1216
			"00000000000000001000000111011010" , -- ADDR 1217
			"00000000000000010001010000110111" , -- ADDR 1218
			"00000000000000001000101010001100" , -- ADDR 1219
			"00000000000000001000000101110000" , -- ADDR 1220
			"00000000000000000101100100111111" , -- ADDR 1221
			"00000000000000001000011001101001" , -- ADDR 1222
			"00000000000000000101010010000001" , -- ADDR 1223
			"00000000000000010011001101111011" , -- ADDR 1224
			"00000000000000001000000111011010" , -- ADDR 1225
			"00000000000000001111011101011101" , -- ADDR 1226
			"00000000000000001010101100110101" , -- ADDR 1227
			"00000000000000001111001111100010" , -- ADDR 1228
			"00000000000000000100001010000101" , -- ADDR 1229
			"00000000000000000101110010011011" , -- ADDR 1230
			"00000000000000000101101000101111" , -- ADDR 1231
			"00000000000000001110000101101010" , -- ADDR 1232
			"00000000000000001110101010110011" , -- ADDR 1233
			"00000000000000001001111001001010" , -- ADDR 1234
			"00000000000000001100101010101100" , -- ADDR 1235
			"00000000000000000111100001010110" , -- ADDR 1236
			"00000000000000000111101000001001" , -- ADDR 1237
			"00000000000000010001000010110110" , -- ADDR 1238
			"00000000000000010010011111011111" , -- ADDR 1239
			"00000000000000000100010001010101" , -- ADDR 1240
			"00000000000000000110001110010111" , -- ADDR 1241
			"00000000000000010111010100100101" , -- ADDR 1242
			"00000000000000001101101100011001" , -- ADDR 1243
			"00000000000000010011001111100000" , -- ADDR 1244
			"00000000000000001110101001101000" , -- ADDR 1245
			"00000000000000000101001001100111" , -- ADDR 1246
			"00000000000000010001110101111010" , -- ADDR 1247
			"00000000000000000011111100011011" , -- ADDR 1248
			"00000000000000001011000000101100" , -- ADDR 1249
			"00000000000000001110010111000110" , -- ADDR 1250
			"00000000000000001110000001101110" , -- ADDR 1251
			"00000000000000000101100111101110" , -- ADDR 1252
			"00000000000000000110101101111010" , -- ADDR 1253
			"00000000000000000111010000100100" , -- ADDR 1254
			"00000000000000000001111101111110" , -- ADDR 1255
			"00000000000000010101001100110001" , -- ADDR 1256
			"00000000000000010011001010011100" , -- ADDR 1257
			"00000000000000001010000101111100" , -- ADDR 1258
			"00000000000000001001100100110001" , -- ADDR 1259
			"00000000000000001100100000011001" , -- ADDR 1260
			"00000000000000001110101001101000" , -- ADDR 1261
			"00000000000000010101011010101111" , -- ADDR 1262
			"00000000000000010100110000001000" , -- ADDR 1263
			"00000000000000000101010010000001" , -- ADDR 1264
			"00000000000000010001011001010101" , -- ADDR 1265
			"00000000000000001111111111101001" , -- ADDR 1266
			"00000000000000001000100100111000" , -- ADDR 1267
			"00000000000000001100011110010000" , -- ADDR 1268
			"00000000000000001001110001011001" , -- ADDR 1269
			"00000000000000000101011101011001" , -- ADDR 1270
			"00000000000000010000101100111011" , -- ADDR 1271
			"00000000000000010000111111000010" , -- ADDR 1272
			"00000000000000001110101001101000" , -- ADDR 1273
			"00000000000000000100011111010001" , -- ADDR 1274
			"00000000000000000111001011100011" , -- ADDR 1275
			"00000000000000000001011011000111" , -- ADDR 1276
			"00000000000000001011111001111101" , -- ADDR 1277
			"00000000000000010011000010100011" , -- ADDR 1278
			"00000000000000010010101000100010" , -- ADDR 1279
			"00000000000000000001000010010011" , -- ADDR 1280
			"00000000000000010001101000101100" , -- ADDR 1281
			"00000000000000001110100100100010" , -- ADDR 1282
			"00000000000000000001100010110101" , -- ADDR 1283
			"00000000000000010000001010001101" , -- ADDR 1284
			"00000000000000001110110110011100" , -- ADDR 1285
			"00000000000000000011100110101101" , -- ADDR 1286
			"00000000000000000101011111001000" , -- ADDR 1287
			"00000000000000001010011100110010" , -- ADDR 1288
			"00000000000000011000100011111011" , -- ADDR 1289
			"00000000000000010001110001100001" , -- ADDR 1290
			"00000000000000010101010011000011" , -- ADDR 1291
			"00000000000000010010011110010000" , -- ADDR 1292
			"00000000000000000011000011110010" , -- ADDR 1293
			"00000000000000010100111101010011" , -- ADDR 1294
			"00000000000000000011101010011000" , -- ADDR 1295
			"00000000000000001110101110001011" , -- ADDR 1296
			"00000000000000001110000001010100" , -- ADDR 1297
			"00000000000000001110101100110000" , -- ADDR 1298
			"00000000000000000110110110100111" , -- ADDR 1299
			"00000000000000000010101011111000" , -- ADDR 1300
			"00000000000000000100110010111111" , -- ADDR 1301
			"00000000000000000010100110000110" , -- ADDR 1302
			"00000000000000010110001010100001" , -- ADDR 1303
			"00000000000000010100100101011011" , -- ADDR 1304
			"00000000000000001100100111001110" , -- ADDR 1305
			"00000000000000001100101110111010" , -- ADDR 1306
			"00000000000000001110100011011111" , -- ADDR 1307
			"00000000000000010001011110100101" , -- ADDR 1308
			"00000000000000010110101101001101" , -- ADDR 1309
			"00000000000000010110101101011110" , -- ADDR 1310
			"00000000000000000010010100001111" , -- ADDR 1311
			"00000000000000001111111110110100" , -- ADDR 1312
			"00000000000000010100000101101000" , -- ADDR 1313
			"00000000000000000110111111011100" , -- ADDR 1314
			"00000000000000001010101010100001" , -- ADDR 1315
			"00000000000000001001011000010011" , -- ADDR 1316
			"00000000000000000110101010110001" , -- ADDR 1317
			"00000000000000010000000101000111" , -- ADDR 1318
			"00000000000000010101001011001001" , -- ADDR 1319
			"00000000000000001100111010010111" , -- ADDR 1320
			"00000000000000001000101100011001" , -- ADDR 1321
			"00000000000000000100110111010101" , -- ADDR 1322
			"00000000000000000100100000000111" , -- ADDR 1323
			"00000000000000001011100001100010" , -- ADDR 1324
			"00000000000000010100001101110001" , -- ADDR 1325
			"00000000000000010010011010111100" , -- ADDR 1326
			"00000000000000000101010010000001" , -- ADDR 1327
			"00000000000000001110011101011100" , -- ADDR 1328
			"00000000000000001100010010110111" , -- ADDR 1329
			"00000000000000000101011001111000" , -- ADDR 1330
			"00000000000000001110101111110111" , -- ADDR 1331
			"00000000000000010001011110010000" , -- ADDR 1332
			"00000000000000000011111011111101" , -- ADDR 1333
			"00000000000000000100011001101100" , -- ADDR 1334
			"00000000000000011000000001101100" , -- ADDR 1335
			"00000000000000001000111010010001" , -- ADDR 1336
			"00000000000000010010111001101101" , -- ADDR 1337
			"00000000000000001010101111101011" , -- ADDR 1338
			"00000000000000001010011011100000" , -- ADDR 1339
			"00000000000000001111100001110000" , -- ADDR 1340
			"00000000000000001000101110010111" , -- ADDR 1341
			"00000000000000001000000000100010" , -- ADDR 1342
			"00000000000000010001110100101111" , -- ADDR 1343
			"00000000000000010000010101011110" , -- ADDR 1344
			"00000000000000000111110100111110" , -- ADDR 1345
			"00000000000000001100101100000011" , -- ADDR 1346
			"00000000000000001101000100011111" , -- ADDR 1347
			"00000000000000000111111011000010" , -- ADDR 1348
			"00000000000000010110011100010100" , -- ADDR 1349
			"00000000000000010011110111110010" , -- ADDR 1350
			"00000000000000001010010010101010" , -- ADDR 1351
			"00000000000000001000100010101010" , -- ADDR 1352
			"00000000000000001101000000111110" , -- ADDR 1353
			"00000000000000001101010100100010" , -- ADDR 1354
			"00000000000000010110001010100001" , -- ADDR 1355
			"00000000000000010100011101100111" , -- ADDR 1356
			"00000000000000001011011010100011" , -- ADDR 1357
			"00000000000000010101101101111011" , -- ADDR 1358
			"00000000000000001011000000101100" , -- ADDR 1359
			"00000000000000001101110010001110" , -- ADDR 1360
			"00000000000000010001011100101110" , -- ADDR 1361
			"00000000000000001101111000110110" , -- ADDR 1362
			"00000000000000001001010010111111" , -- ADDR 1363
			"00000000000000010100010000111110" , -- ADDR 1364
			"00000000000000001011100010100001" , -- ADDR 1365
			"00000000000000010011011011000011" , -- ADDR 1366
			"00000000000000000001110000101011" , -- ADDR 1367
			"00000000000000001100111100001000" , -- ADDR 1368
			"00000000000000000110000111100100" , -- ADDR 1369
			"00000000000000001111101100011001" , -- ADDR 1370
			"00000000000000010100001000011110" , -- ADDR 1371
			"00000000000000010101100110001011" , -- ADDR 1372
			"00000000000000000101001100001100" , -- ADDR 1373
			"00000000000000010111011000011011" , -- ADDR 1374
			"00000000000000010011110001100010" , -- ADDR 1375
			"00000000000000000101100111101110" , -- ADDR 1376
			"00000000000000010100100011001100" , -- ADDR 1377
			"00000000000000001101111010110001" , -- ADDR 1378
			"00000000000000001000001011110110" , -- ADDR 1379
			"00000000000000001010000000101000" , -- ADDR 1380
			"00000000000000010011111011001111" , -- ADDR 1381
			"00000000000000000101110111010101" , -- ADDR 1382
			"00000000000000010001011000001000" , -- ADDR 1383
			"00000000000000011011011000100001" , -- ADDR 1384
			"00000000000000001100000001100110" , -- ADDR 1385
			"00000000000000011010111100001001" , -- ADDR 1386
			"00000000000000010001000100100001" , -- ADDR 1387
			"00000000000000001011111110010001" , -- ADDR 1388
			"00000000000000001001111101110001" , -- ADDR 1389
			"00000000000000011100111001000111" , -- ADDR 1390
			"00000000000000011010101111110010" , -- ADDR 1391
			"00000000000000010100111111000111" , -- ADDR 1392
			"00000000000000011000100001100001" , -- ADDR 1393
			"00000000000000000010101110101100" , -- ADDR 1394
			"00000000000000000100001100110101" , -- ADDR 1395
			"00000000000000001101110100011100" , -- ADDR 1396
			"00000000000000001111100000010010" , -- ADDR 1397
			"00000000000000001011000110101110" , -- ADDR 1398
			"00000000000000001011011111100010" , -- ADDR 1399
			"00000000000000000001111010000010" , -- ADDR 1400
			"00000000000000000100101100100011" , -- ADDR 1401
			"00000000000000010110101011110010" , -- ADDR 1402
			"00000000000000001110011010000000" , -- ADDR 1403
			"00000000000000010100100000100110" , -- ADDR 1404
			"00000000000000010010101010111111" , -- ADDR 1405
			"00000000000000010001001111001101" , -- ADDR 1406
			"00000000000000001111101000001000" , -- ADDR 1407
			"00000000000000010010001001011010" , -- ADDR 1408
			"00000000000000001011100001000010" , -- ADDR 1409
			"00000000000000010110011101100101" , -- ADDR 1410
			"00000000000000010000010011000001" , -- ADDR 1411
			"00000000000000010111111010011000" , -- ADDR 1412
			"00000000000000010100110001100000" , -- ADDR 1413
			"00000000000000011000101101110101" , -- ADDR 1414
			"00000000000000001101111000011011" , -- ADDR 1415
			"00000000000000000100010110001100" , -- ADDR 1416
			"00000000000000001001000010010110" , -- ADDR 1417
			"00000000000000010111011000100000" , -- ADDR 1418
			"00000000000000010110011110010001" , -- ADDR 1419
			"00000000000000010010010000111101" , -- ADDR 1420
			"00000000000000010101111110101100" , -- ADDR 1421
			"00000000000000001110101011100101" , -- ADDR 1422
			"00000000000000001010100110011001" , -- ADDR 1423
			"00000000000000011010110000100100" , -- ADDR 1424
			"00000000000000011100010110000111" , -- ADDR 1425
			"00000000000000001110000101101010" , -- ADDR 1426
			"00000000000000000010101110101100" , -- ADDR 1427
			"00000000000000010010101011110011" , -- ADDR 1428
			"00000000000000001000101000001101" , -- ADDR 1429
			"00000000000000010001001000100010" , -- ADDR 1430
			"00000000000000000100001100110101" , -- ADDR 1431
			"00000000000000010010101011111010" , -- ADDR 1432
			"00000000000000001111110111101000" , -- ADDR 1433
			"00000000000000010000101101110101" , -- ADDR 1434
			"00000000000000010100010111101001" , -- ADDR 1435
			"00000000000000010010100000011010" , -- ADDR 1436
			"00000000000000001111101010000101" , -- ADDR 1437
			"00000000000000010011010010011110" , -- ADDR 1438
			"00000000000000010000010110111000" , -- ADDR 1439
			"00000000000000001001011010111100" , -- ADDR 1440
			"00000000000000000111010100110000" , -- ADDR 1441
			"00000000000000001011000111100101" , -- ADDR 1442
			"00000000000000001000100010111000" , -- ADDR 1443
			"00000000000000010010010110011110" , -- ADDR 1444
			"00000000000000001111011101110100" , -- ADDR 1445
			"00000000000000010001110100101111" , -- ADDR 1446
			"00000000000000010111010100100101" , -- ADDR 1447
			"00000000000000000010010100001111" , -- ADDR 1448
			"00000000000000010010000100101011" , -- ADDR 1449
			"00000000000000010100101110100100" , -- ADDR 1450
			"00000000000000010000100101100101" , -- ADDR 1451
			"00000000000000001101010101110100" , -- ADDR 1452
			"00000000000000010100110110110100" , -- ADDR 1453
			"00000000000000000011110011000100" , -- ADDR 1454
			"00000000000000010110000100111011" , -- ADDR 1455
			"00000000000000001010010001000000" , -- ADDR 1456
			"00000000000000010010010011000011" , -- ADDR 1457
			"00000000000000001110001111000110" , -- ADDR 1458
			"00000000000000010001011110111010" , -- ADDR 1459
			"00000000000000010001000111100010" , -- ADDR 1460
			"00000000000000010101000100111011" , -- ADDR 1461
			"00000000000000001100110110000100" , -- ADDR 1462
			"00000000000000011011101000010100" , -- ADDR 1463
			"00000000000000010111001001111111" , -- ADDR 1464
			"00000000000000001100011000000111" , -- ADDR 1465
			"00000000000000010110011010100010" , -- ADDR 1466
			"00000000000000001001100001100101" , -- ADDR 1467
			"00000000000000010000101000010110" , -- ADDR 1468
			"00000000000000010010100100011011" , -- ADDR 1469
			"00000000000000001011100001000010" , -- ADDR 1470
			"00000000000000010111110101010001" , -- ADDR 1471
			"00000000000000000110010001101110" , -- ADDR 1472
			"00000000000000010111000101110010" , -- ADDR 1473
			"00000000000000001011011110100011" , -- ADDR 1474
			"00000000000000001011011111100010" , -- ADDR 1475
			"00000000000000001000010101010100" , -- ADDR 1476
			"00000000000000011000100110011111" , -- ADDR 1477
			"00000000000000010111110000011101" , -- ADDR 1478
			"00000000000000010010100101111110" , -- ADDR 1479
			"00000000000000010100101110101010" , -- ADDR 1480
			"00000000000000000101111001100110" , -- ADDR 1481
			"00000000000000000011010010001110" , -- ADDR 1482
			"00000000000000001001001100001011" , -- ADDR 1483
			"00000000000000001010011010001110" , -- ADDR 1484
			"00000000000000000110110010001001" , -- ADDR 1485
			"00000000000000000101110011011010" , -- ADDR 1486
			"00000000000000000100100000000111" , -- ADDR 1487
			"00000000000000000001100100000011" , -- ADDR 1488
			"00000000000000010011110001100010" , -- ADDR 1489
			"00000000000000001111011010110111" , -- ADDR 1490
			"00000000000000001110101001100000" , -- ADDR 1491
			"00000000000000010000100100111001" , -- ADDR 1492
			"00000000000000010000011001110010" , -- ADDR 1493
			"00000000000000001101100010010100" , -- ADDR 1494
			"00000000000000001110101000011101" , -- ADDR 1495
			"00000000000000001100001111110000" , -- ADDR 1496
			"00000000000000010000100110111101" , -- ADDR 1497
			"00000000000000010000001110111011" , -- ADDR 1498
			"00000000000000010011000010100011" , -- ADDR 1499
			"00000000000000010010010110110010" , -- ADDR 1500
			"00000000000000010100100011101010" , -- ADDR 1501
			"00000000000000001100011101000010" , -- ADDR 1502
			"00000000000000000100011111010001" , -- ADDR 1503
			"00000000000000001010101100110101" , -- ADDR 1504
			"00000000000000010011000110100011" , -- ADDR 1505
			"00000000000000010110110011010000" , -- ADDR 1506
			"00000000000000010010000110100100" , -- ADDR 1507
			"00000000000000010001110001100001" , -- ADDR 1508
			"00000000000000001111001101011010" , -- ADDR 1509
			"00000000000000000101000001101111" , -- ADDR 1510
			"00000000000000010110110100100101" , -- ADDR 1511
			"00000000000000011000100101011111" , -- ADDR 1512
			"00000000000000010011110001101110" , -- ADDR 1513
			"00000000000000000101111001100110" , -- ADDR 1514
			"00000000000000010010010110011110" , -- ADDR 1515
			"00000000000000000011110010100100" , -- ADDR 1516
			"00000000000000010001010010010011" , -- ADDR 1517
			"00000000000000001110001111000110" , -- ADDR 1518
			"00000000000000010010010110110010" , -- ADDR 1519
			"00000000000000010101001000110011" , -- ADDR 1520
			"00000000000000010010011111111001" , -- ADDR 1521
			"00000000000000010000100110111101" , -- ADDR 1522
			"00000000000000010000111010001100" , -- ADDR 1523
			"00000000000000001101111110000011" , -- ADDR 1524
			"00000000000000001000010010110011" , -- ADDR 1525
			"00000000000000000110100100101110" , -- ADDR 1526
			"00000000000000001001011010111100" , -- ADDR 1527
			"00000000000000000110001110010111" , -- ADDR 1528
			"00000000000000001111110111101000" , -- ADDR 1529
			"00000000000000001100110110000100" , -- ADDR 1530
			"00000000000000010010001011100001" , -- ADDR 1531
			"00000000000000010101111110010000" , -- ADDR 1532
			"00000000000000000011010100100001" , -- ADDR 1533
			"00000000000000010001101101110000" , -- ADDR 1534
			"00000000000000010011111100011000" , -- ADDR 1535
			"00000000000000001111110100101111" , -- ADDR 1536
			"00000000000000001101001111010111" , -- ADDR 1537
			"00000000000000010011010011100100" , -- ADDR 1538
			"00000000000000000101010101010000" , -- ADDR 1539
			"00000000000000010101000011111011" , -- ADDR 1540
			"00000000000000001011110101111100" , -- ADDR 1541
			"00000000000000010010010001011111" , -- ADDR 1542
			"00000000000000001111011010010111" , -- ADDR 1543
			"00000000000000010000011001101011" , -- ADDR 1544
			"00000000000000001110110011111111" , -- ADDR 1545
			"00000000000000010011001111000111" , -- ADDR 1546
			"00000000000000001101111011001011" , -- ADDR 1547
			"00000000000000011010111101010110" , -- ADDR 1548
			"00000000000000010110010100101111" , -- ADDR 1549
			"00000000000000001101001101000011" , -- ADDR 1550
			"00000000000000010101001010011011" , -- ADDR 1551
			"00000000000000000111001110101110" , -- ADDR 1552
			"00000000000000010001111000011110" , -- ADDR 1553
			"00000000000000010011110110010110" , -- ADDR 1554
			"00000000000000010110111010100110" , -- ADDR 1555
			"00000000000000000001110000101011" , -- ADDR 1556
			"00000000000000010000001010001101" , -- ADDR 1557
			"00000000000000010001000100000101" , -- ADDR 1558
			"00000000000000010001100110111101" , -- ADDR 1559
			"00000000000000000100100101100100" , -- ADDR 1560
			"00000000000000000010111100110011" , -- ADDR 1561
			"00000000000000000111110011010001" , -- ADDR 1562
			"00000000000000000011010000011110" , -- ADDR 1563
			"00000000000000011001000010111111" , -- ADDR 1564
			"00000000000000010111010101110011" , -- ADDR 1565
			"00000000000000001110110111111110" , -- ADDR 1566
			"00000000000000001110101000000100" , -- ADDR 1567
			"00000000000000010001000011001100" , -- ADDR 1568
			"00000000000000010011100111000100" , -- ADDR 1569
			"00000000000000011001100000100100" , -- ADDR 1570
			"00000000000000011001010010100010" , -- ADDR 1571
			"00000000000000000101010110101100" , -- ADDR 1572
			"00000000000000010011000000001001" , -- ADDR 1573
			"00000000000000010100111101010011" , -- ADDR 1574
			"00000000000000001010000010111010" , -- ADDR 1575
			"00000000000000001101101010100101" , -- ADDR 1576
			"00000000000000001100011001110100" , -- ADDR 1577
			"00000000000000001001010001111101" , -- ADDR 1578
			"00000000000000010011001000110110" , -- ADDR 1579
			"00000000000000010101110010110101" , -- ADDR 1580
			"00000000000000001111111001111010" , -- ADDR 1581
			"00000000000000001000101110010111" , -- ADDR 1582
			"00000000000000000111111000110111" , -- ADDR 1583
			"00000000000000000100011101001000" , -- ADDR 1584
			"00000000000000001110100011111001" , -- ADDR 1585
			"00000000000000010111000010011110" , -- ADDR 1586
			"00000000000000010101011101110000" , -- ADDR 1587
			"00000000000000000101110111010101" , -- ADDR 1588
			"00000000000000010000111010001100" , -- ADDR 1589
			"00000000000000001111001011011001" , -- ADDR 1590
			"00000000000000000110101010011111" , -- ADDR 1591
			"00000000000000010001110001100001" , -- ADDR 1592
			"00000000000000010011101110001001" , -- ADDR 1593
			"00000000000000000010010011011010" , -- ADDR 1594
			"00000000000000000001011101110000" , -- ADDR 1595
			"00000000000000010101110001100001" , -- ADDR 1596
			"00000000000000000111100001010110" , -- ADDR 1597
			"00000000000000001111010011011010" , -- ADDR 1598
			"00000000000000001011111010111010" , -- ADDR 1599
			"00000000000000010110011111101000" , -- ADDR 1600
			"00000000000000010111100111101011" , -- ADDR 1601
			"00000000000000010011100110110010" , -- ADDR 1602
			"00000000000000010011101010001011" , -- ADDR 1603
			"00000000000000001100000111110001" , -- ADDR 1604
			"00000000000000001001010010111111" , -- ADDR 1605
			"00000000000000001000100011000110" , -- ADDR 1606
			"00000000000000001000010010100100" , -- ADDR 1607
			"00000000000000000111110011010001" , -- ADDR 1608
			"00000000000000000011101111000001" , -- ADDR 1609
			"00000000000000001010110001110011" , -- ADDR 1610
			"00000000000000000111010101110011" , -- ADDR 1611
			"00000000000000010100000010000111" , -- ADDR 1612
			"00000000000000010011110101000000" , -- ADDR 1613
			"00000000000000001000101010110111" , -- ADDR 1614
			"00000000000000010010001001011010" , -- ADDR 1615
			"00000000000000010011010001001100" , -- ADDR 1616
			"00000000000000001111100001110000" , -- ADDR 1617
			"00000000000000001110101001101000" , -- ADDR 1618
			"00000000000000010000110010100000" , -- ADDR 1619
			"00000000000000001010100010110010" , -- ADDR 1620
			"00000000000000010011110001101110" , -- ADDR 1621
			"00000000000000010000001101000010" , -- ADDR 1622
			"00000000000000010011010111001110" , -- ADDR 1623
			"00000000000000010010111010110100" , -- ADDR 1624
			"00000000000000001111010010111010" , -- ADDR 1625
			"00000000000000001010010111110101" , -- ADDR 1626
			"00000000000000001111111100010011" , -- ADDR 1627
			"00000000000000010001011000000001" , -- ADDR 1628
			"00000000000000011010001101011011" , -- ADDR 1629
			"00000000000000010101011001110000" , -- ADDR 1630
			"00000000000000010000010011001001" , -- ADDR 1631
			"00000000000000010011010011010001" , -- ADDR 1632
			"00000000000000000100010000111000" , -- ADDR 1633
			"00000000000000010101011000101100" , -- ADDR 1634
			"00000000000000010111010100010101" , -- ADDR 1635
			"00000000000000001110110011111111" , -- ADDR 1636
			"00000000000000010001001001011011" , -- ADDR 1637
			"00000000000000010001010110010111" , -- ADDR 1638
			"00000000000000000011001101100001" , -- ADDR 1639
			"00000000000000000100100010101001" , -- ADDR 1640
			"00000000000000001000011000111110" , -- ADDR 1641
			"00000000000000000010011010101011" , -- ADDR 1642
			"00000000000000011000101100111010" , -- ADDR 1643
			"00000000000000010110110101000101" , -- ADDR 1644
			"00000000000000001101111111011010" , -- ADDR 1645
			"00000000000000001101100001000010" , -- ADDR 1646
			"00000000000000010000010100100011" , -- ADDR 1647
			"00000000000000010010100101111110" , -- ADDR 1648
			"00000000000000011001000010111111" , -- ADDR 1649
			"00000000000000011000100101010000" , -- ADDR 1650
			"00000000000000000101111001111011" , -- ADDR 1651
			"00000000000000010011011111000100" , -- ADDR 1652
			"00000000000000010011011000101100" , -- ADDR 1653
			"00000000000000001010011011100000" , -- ADDR 1654
			"00000000000000001110001110001001" , -- ADDR 1655
			"00000000000000001100011100111000" , -- ADDR 1656
			"00000000000000001000110011100101" , -- ADDR 1657
			"00000000000000010011010101100010" , -- ADDR 1658
			"00000000000000010100001010000101" , -- ADDR 1659
			"00000000000000010000011110001101" , -- ADDR 1660
			"00000000000000000111000010111110" , -- ADDR 1661
			"00000000000000001000011011011101" , -- ADDR 1662
			"00000000000000000010111100001010" , -- ADDR 1663
			"00000000000000001110101000100110" , -- ADDR 1664
			"00000000000000010110100111011010" , -- ADDR 1665
			"00000000000000010101100010000001" , -- ADDR 1666
			"00000000000000000100011101001000" , -- ADDR 1667
			"00000000000000010010000011111100" , -- ADDR 1668
			"00000000000000001111111011111100" , -- ADDR 1669
			"00000000000000000101011111001000" , -- ADDR 1670
			"00000000000000010010001111100110" , -- ADDR 1671
			"00000000000000010010110001111010" , -- ADDR 1672
			"00000000000000000000100010111100" , -- ADDR 1673
			"00000000000000000001100010110101" , -- ADDR 1674
			"00000000000000001110100001011001" , -- ADDR 1675
			"00000000000000001011110100000000" , -- ADDR 1676
			"00000000000000001111001001010000" , -- ADDR 1677
			"00000000000000010001011001010101" , -- ADDR 1678
			"00000000000000001110101111111111" , -- ADDR 1679
			"00000000000000001100111100101110" , -- ADDR 1680
			"00000000000000010000000001010100" , -- ADDR 1681
			"00000000000000001101001010101111" , -- ADDR 1682
			"00000000000000000101001111011111" , -- ADDR 1683
			"00000000000000000011001000000110" , -- ADDR 1684
			"00000000000000000111001011110100" , -- ADDR 1685
			"00000000000000000101101011011011" , -- ADDR 1686
			"00000000000000001111010101100001" , -- ADDR 1687
			"00000000000000001100111111101010" , -- ADDR 1688
			"00000000000000001110011000111101" , -- ADDR 1689
			"00000000000000010011001000110110" , -- ADDR 1690
			"00000000000000000110001110010111" , -- ADDR 1691
			"00000000000000001110000101011001" , -- ADDR 1692
			"00000000000000010000100100101010" , -- ADDR 1693
			"00000000000000001100011011100000" , -- ADDR 1694
			"00000000000000001001011111111110" , -- ADDR 1695
			"00000000000000010000101110111110" , -- ADDR 1696
			"00000000000000000111111110001010" , -- ADDR 1697
			"00000000000000010001111000011110" , -- ADDR 1698
			"00000000000000001000101111000001" , -- ADDR 1699
			"00000000000000001110100001110010" , -- ADDR 1700
			"00000000000000001011111000010110" , -- ADDR 1701
			"00000000000000001101010010000110" , -- ADDR 1702
			"00000000000000001101110000000001" , -- ADDR 1703
			"00000000000000010001000111001101" , -- ADDR 1704
			"00000000000000001010010110111010" , -- ADDR 1705
			"00000000000000010111100001001101" , -- ADDR 1706
			"00000000000000010010111111100011" , -- ADDR 1707
			"00000000000000001001100001100101" , -- ADDR 1708
			"00000000000000010010001110000010" , -- ADDR 1709
			"00000000000000000110011111001011" , -- ADDR 1710
			"00000000000000001110010111101000" , -- ADDR 1711
			"00000000000000010000010101011110" , -- ADDR 1712
			"00000000000000000011011001000100" , -- ADDR 1713
			"00000000000000010011110100000010" , -- ADDR 1714
			"00000000000000001111101101111110" , -- ADDR 1715
			"00000000000000001001101010101110" , -- ADDR 1716
			"00000000000000001110110110100100" , -- ADDR 1717
			"00000000000000001001010000111011" , -- ADDR 1718
			"00000000000000001001000010001000" , -- ADDR 1719
			"00000000000000001001010001111101" , -- ADDR 1720
			"00000000000000001011011110100011" , -- ADDR 1721
			"00000000000000000111111100101110" , -- ADDR 1722
			"00000000000000001011111100010110" , -- ADDR 1723
			"00000000000000001010011100000011" , -- ADDR 1724
			"00000000000000001100010001001001" , -- ADDR 1725
			"00000000000000001011110100011111" , -- ADDR 1726
			"00000000000000000100101100001001" , -- ADDR 1727
			"00000000000000010100011100110010" , -- ADDR 1728
			"00000000000000000111010000000010" , -- ADDR 1729
			"00000000000000000101010001010011" , -- ADDR 1730
			"00000000000000000100101100100011" , -- ADDR 1731
			"00000000000000001001000000001110" , -- ADDR 1732
			"00000000000000000010011100010000" , -- ADDR 1733
			"00000000000000010110010111000010" , -- ADDR 1734
			"00000000000000000100101111011000" , -- ADDR 1735
			"00000000000000010000111000111101" , -- ADDR 1736
			"00000000000000001001011111110001" , -- ADDR 1737
			"00000000000000001111110000000010" , -- ADDR 1738
			"00000000000000000010100000111000" , -- ADDR 1739
			"00000000000000001000000101110000" , -- ADDR 1740
			"00000000000000000100011001101100" , -- ADDR 1741
			"00000000000000001110110111001101" , -- ADDR 1742
			"00000000000000001011010011110101" , -- ADDR 1743
			"00000000000000000110101000011110" , -- ADDR 1744
			"00000000000000001101100000010101" , -- ADDR 1745
			"00000000000000000100000000010001" , -- ADDR 1746
			"00000000000000001011001000100111" , -- ADDR 1747
			"00000000000000010001001001000110" , -- ADDR 1748
			"00000000000000010010010011000011" , -- ADDR 1749
			"00000000000000010011101001000111" , -- ADDR 1750
			"00000000000000010000110011010011" , -- ADDR 1751
			"00000000000000001011000001111001" , -- ADDR 1752
			"00000000000000001110111100100101" , -- ADDR 1753
			"00000000000000000111011110010010" , -- ADDR 1754
			"00000000000000000110010101101010" , -- ADDR 1755
			"00000000000000000110101101000011" , -- ADDR 1756
			"00000000000000001000111101000010" , -- ADDR 1757
			"00000000000000000100110100001011" , -- ADDR 1758
			"00000000000000001000101000011011" , -- ADDR 1759
			"00000000000000001000001100000101" , -- ADDR 1760
			"00000000000000001001010010100101" , -- ADDR 1761
			"00000000000000001100101111101010" , -- ADDR 1762
			"00000000000000000111111100101110" , -- ADDR 1763
			"00000000000000010001011110100101" , -- ADDR 1764
			"00000000000000001000110000000111" , -- ADDR 1765
			"00000000000000001000000100100101" , -- ADDR 1766
			"00000000000000000101101011011011" , -- ADDR 1767
			"00000000000000001000100110011100" , -- ADDR 1768
			"00000000000000000101000101001001" , -- ADDR 1769
			"00000000000000010011011011110101" , -- ADDR 1770
			"00000000000000001000000001111110" , -- ADDR 1771
			"00000000000000001111101100100000" , -- ADDR 1772
			"00000000000000001010110100000110" , -- ADDR 1773
			"00000000000000001111011100110101" , -- ADDR 1774
			"00000000000000000100001011011101" , -- ADDR 1775
			"00000000000000000101101011011011" , -- ADDR 1776
			"00000000000000000101011001001011" , -- ADDR 1777
			"00000000000000001110010011100000" , -- ADDR 1778
			"00000000000000001110100101111111" , -- ADDR 1779
			"00000000000000001001110101000110" , -- ADDR 1780
			"00000000000000001100111000100101" , -- ADDR 1781
			"00000000000000000111011000011000" , -- ADDR 1782
			"00000000000000000111110010010010" , -- ADDR 1783
			"00000000000000010001001111001101" , -- ADDR 1784
			"00000000000000010010101011000101" , -- ADDR 1785
			"00000000000000000111100010010111" , -- ADDR 1786
			"00000000000000001011011111111000" , -- ADDR 1787
			"00000000000000000101000010001000" , -- ADDR 1788
			"00000000000000011010110011110001" , -- ADDR 1789
			"00000000000000011000101101110101" , -- ADDR 1790
			"00000000000000001111011010010111" , -- ADDR 1791
			"00000000000000001110011111100011" , -- ADDR 1792
			"00000000000000010001111101010001" , -- ADDR 1793
			"00000000000000010011101001000111" , -- ADDR 1794
			"00000000000000011010111111000111" , -- ADDR 1795
			"00000000000000011010001000110000" , -- ADDR 1796
			"00000000000000001001000010010110" , -- ADDR 1797
			"00000000000000010110011101010000" , -- ADDR 1798
			"00000000000000010010110101101010" , -- ADDR 1799
			"00000000000000001101011010000110" , -- ADDR 1800
			"00000000000000010001010000110111" , -- ADDR 1801
			"00000000000000001111001001010000" , -- ADDR 1802
			"00000000000000001011000011011101" , -- ADDR 1803
			"00000000000000010110000101101101" , -- ADDR 1804
			"00000000000000010011010011010001" , -- ADDR 1805
			"00000000000000010011100000100010" , -- ADDR 1806
			"00000000000000000110100000111011" , -- ADDR 1807
			"00000000000000001011100001000010" , -- ADDR 1808
			"00000000000000000100001100110101" , -- ADDR 1809
			"00000000000000010001010100011001" , -- ADDR 1810
			"00000000000000011000101000100000" , -- ADDR 1811
			"00000000000000011000001001010011" , -- ADDR 1812
			"00000000000000000101100001100011" , -- ADDR 1813
			"00000000000000010101010001011100" , -- ADDR 1814
			"00000000000000010011000100010110" , -- ADDR 1815
			"00000000000000000110111010100000" , -- ADDR 1816
			"00000000000000010101001101100101" , -- ADDR 1817
			"00000000000000010011111110110001" , -- ADDR 1818
			"00000000000000000010111011100000" , -- ADDR 1819
			"00000000000000000011010100100001" , -- ADDR 1820
			"00000000000000000110000100000111" , -- ADDR 1821
			"00000000000000000100110011110010" , -- ADDR 1822
			"00000000000000011000010001001011" , -- ADDR 1823
			"00000000000000010110110111010000" , -- ADDR 1824
			"00000000000000001111001110100010" , -- ADDR 1825
			"00000000000000001111011010010111" , -- ADDR 1826
			"00000000000000010001000100000101" , -- ADDR 1827
			"00000000000000010100000111001001" , -- ADDR 1828
			"00000000000000011000111011000011" , -- ADDR 1829
			"00000000000000011001001000101100" , -- ADDR 1830
			"00000000000000000100000100000011" , -- ADDR 1831
			"00000000000000010001000010001011" , -- ADDR 1832
			"00000000000000010110101011011100" , -- ADDR 1833
			"00000000000000001000011110011001" , -- ADDR 1834
			"00000000000000001011101100001101" , -- ADDR 1835
			"00000000000000001011010000010010" , -- ADDR 1836
			"00000000000000001001001100001011" , -- ADDR 1837
			"00000000000000010001100101000111" , -- ADDR 1838
			"00000000000000010111101100111010" , -- ADDR 1839
			"00000000000000001101110111011110" , -- ADDR 1840
			"00000000000000001010111011101001" , -- ADDR 1841
			"00000000000000000110001110010111" , -- ADDR 1842
			"00000000000000000110100100101110" , -- ADDR 1843
			"00000000000000001101010010110100" , -- ADDR 1844
			"00000000000000010110011010100010" , -- ADDR 1845
			"00000000000000010100000100101011" , -- ADDR 1846
			"00000000000000000111101010011001" , -- ADDR 1847
			"00000000000000001110001010011001" , -- ADDR 1848
			"00000000000000001100111001001011" , -- ADDR 1849
			"00000000000000000111111111110101" , -- ADDR 1850
			"00000000000000001111110101110101" , -- ADDR 1851
			"00000000000000010100000100110001" , -- ADDR 1852
			"00000000000000000101000010001000" , -- ADDR 1853
			"00000000000000000100010100111000" , -- ADDR 1854
			"00000000000000000110100111000010" , -- ADDR 1855
			"00000000000000010010011011010000" , -- ADDR 1856
			"00000000000000010001010001110110" , -- ADDR 1857
			"00000000000000001011000101010110" , -- ADDR 1858
			"00000000000000001100000010111000" , -- ADDR 1859
			"00000000000000001100001111110000" , -- ADDR 1860
			"00000000000000001111111001100011" , -- ADDR 1861
			"00000000000000010011001101111011" , -- ADDR 1862
			"00000000000000010011110110101000" , -- ADDR 1863
			"00000000000000000010011111010110" , -- ADDR 1864
			"00000000000000001011001100111000" , -- ADDR 1865
			"00000000000000010100110001100000" , -- ADDR 1866
			"00000000000000000010011010101011" , -- ADDR 1867
			"00000000000000000101110111101010" , -- ADDR 1868
			"00000000000000000101010111000010" , -- ADDR 1869
			"00000000000000000101010000100101" , -- ADDR 1870
			"00000000000000001011100001100010" , -- ADDR 1871
			"00000000000000010110001101011101" , -- ADDR 1872
			"00000000000000001000000111011010" , -- ADDR 1873
			"00000000000000001011011110100011" , -- ADDR 1874
			"00000000000000000000001111101000" , -- ADDR 1875
			"00000000000000001000001111000110" , -- ADDR 1876
			"00000000000000000111010010001001" , -- ADDR 1877
			"00000000000000010000101101001001" , -- ADDR 1878
			"00000000000000001110000000101001" , -- ADDR 1879
			"00000000000000001000001101001111" , -- ADDR 1880
			"00000000000000001010011000110000" , -- ADDR 1881
			"00000000000000000111100100101000" , -- ADDR 1882
			"00000000000000000111011101000001" , -- ADDR 1883
			"00000000000000001001111110010101" , -- ADDR 1884
			"00000000000000001111101000000000" , -- ADDR 1885
			"00000000000000001000100100111000" , -- ADDR 1886
			"00000000000000001001001100001011" , -- ADDR 1887
			"00000000000000010110010010010101" , -- ADDR 1888
			"00000000000000010100011010101110" , -- ADDR 1889
			"00000000000000001011101011101110" , -- ADDR 1890
			"00000000000000001011010111101101" , -- ADDR 1891
			"00000000000000001101111100110100" , -- ADDR 1892
			"00000000000000010000010111111011" , -- ADDR 1893
			"00000000000000010110101000011010" , -- ADDR 1894
			"00000000000000010110001101011101" , -- ADDR 1895
			"00000000000000000100010000111000" , -- ADDR 1896
			"00000000000000010001011011011010" , -- ADDR 1897
			"00000000000000010001111101001010" , -- ADDR 1898
			"00000000000000001000011000111110" , -- ADDR 1899
			"00000000000000001100010001001001" , -- ADDR 1900
			"00000000000000001010001010011101" , -- ADDR 1901
			"00000000000000000110011000111101" , -- ADDR 1902
			"00000000000000010001000101110111" , -- ADDR 1903
			"00000000000000010010111010110100" , -- ADDR 1904
			"00000000000000001110100000010110" , -- ADDR 1905
			"00000000000000000110001010010111" , -- ADDR 1906
			"00000000000000000110100110001011" , -- ADDR 1907
			"00000000000000000001111010000010" , -- ADDR 1908
			"00000000000000001100010110000111" , -- ADDR 1909
			"00000000000000010100001100101111" , -- ADDR 1910
			"00000000000000010011001101111011" , -- ADDR 1911
			"00000000000000000010110110111001" , -- ADDR 1912
			"00000000000000010000110001001000" , -- ADDR 1913
			"00000000000000001110001010011001" , -- ADDR 1914
			"00000000000000000011011011010100" , -- ADDR 1915
			"00000000000000010000001011101111" , -- ADDR 1916
			"00000000000000010000100000101000" , -- ADDR 1917
			"00000000000000000010010011011010" , -- ADDR 1918
			"00000000000000000011110111000011" , -- ADDR 1919
			"00000000000000000010111100001010" , -- ADDR 1920
			"00000000000000001100001001101001" , -- ADDR 1921
			"00000000000000001110000011011111" , -- ADDR 1922
			"00000000000000001001011011100010" , -- ADDR 1923
			"00000000000000001010101111101011" , -- ADDR 1924
			"00000000000000000001110000101011" , -- ADDR 1925
			"00000000000000000101011000000111" , -- ADDR 1926
			"00000000000000010100001101110001" , -- ADDR 1927
			"00000000000000001011101111011110" , -- ADDR 1928
			"00000000000000010100001010110000" , -- ADDR 1929
			"00000000000000010000000101000111" , -- ADDR 1930
			"00000000000000001110100001011001" , -- ADDR 1931
			"00000000000000001101000100011111" , -- ADDR 1932
			"00000000000000001111111001011011" , -- ADDR 1933
			"00000000000000001000110011011000" , -- ADDR 1934
			"00000000000000010110001010101100" , -- ADDR 1935
			"00000000000000001101100100011011" , -- ADDR 1936
			"00000000000000010110001010100001" , -- ADDR 1937
			"00000000000000010010001110000010" , -- ADDR 1938
			"00000000000000010110100111001001" , -- ADDR 1939
			"00000000000000001011001111110001" , -- ADDR 1940
			"00000000000000000010010100001111" , -- ADDR 1941
			"00000000000000000110011000111101" , -- ADDR 1942
			"00000000000000010101010101111011" , -- ADDR 1943
			"00000000000000010011110001101110" , -- ADDR 1944
			"00000000000000001111100010011000" , -- ADDR 1945
			"00000000000000010011111011001001" , -- ADDR 1946
			"00000000000000001011111110010001" , -- ADDR 1947
			"00000000000000001001110001000000" , -- ADDR 1948
			"00000000000000011000100011011000" , -- ADDR 1949
			"00000000000000011010000100010111" , -- ADDR 1950
			"00000000000000001001101000010110" , -- ADDR 1951
			"00000000000000001011011000010111" , -- ADDR 1952
			"00000000000000000110111010001110" , -- ADDR 1953
			"00000000000000000111110100000000" , -- ADDR 1954
			"00000000000000000010010011011010" , -- ADDR 1955
			"00000000000000000011011001101000" , -- ADDR 1956
			"00000000000000010010110011100010" , -- ADDR 1957
			"00000000000000001100100000101101" , -- ADDR 1958
			"00000000000000010001001110110000" , -- ADDR 1959
			"00000000000000001111000011110101" , -- ADDR 1960
			"00000000000000001110001101100111" , -- ADDR 1961
			"00000000000000001011111110010001" , -- ADDR 1962
			"00000000000000001110000100011100" , -- ADDR 1963
			"00000000000000001001010110111000" , -- ADDR 1964
			"00000000000000010011001110110100" , -- ADDR 1965
			"00000000000000001101101101001111" , -- ADDR 1966
			"00000000000000010011101110001001" , -- ADDR 1967
			"00000000000000010001000011100001" , -- ADDR 1968
			"00000000000000010100100011001100" , -- ADDR 1969
			"00000000000000001010011111001001" , -- ADDR 1970
			"00000000000000000001001110001000" , -- ADDR 1971
			"00000000000000000111100010100111" , -- ADDR 1972
			"00000000000000010011001100110101" , -- ADDR 1973
			"00000000000000010100001100101111" , -- ADDR 1974
			"00000000000000001111101001000110" , -- ADDR 1975
			"00000000000000010001110011010110" , -- ADDR 1976
			"00000000000000001100011100101110" , -- ADDR 1977
			"00000000000000000110110101110010" , -- ADDR 1978
			"00000000000000010110101000011010" , -- ADDR 1979
			"00000000000000011000010000011110" , -- ADDR 1980
			"00000000000000000010010000000100" , -- ADDR 1981
			"00000000000000000010101110101100" , -- ADDR 1982
			"00000000000000000100111010000100" , -- ADDR 1983
			"00000000000000001011111011101101" , -- ADDR 1984
			"00000000000000001010101110011100" , -- ADDR 1985
			"00000000000000001011100001000010" , -- ADDR 1986
			"00000000000000001101111001101011" , -- ADDR 1987
			"00000000000000001011010010010100" , -- ADDR 1988
			"00000000000000001001110011100010" , -- ADDR 1989
			"00000000000000001011101010111010" , -- ADDR 1990
			"00000000000000000111100101011000" , -- ADDR 1991
			"00000000000000000110000111111000" , -- ADDR 1992
			"00000000000000001011100001000010" , -- ADDR 1993
			"00000000000000001101001001000000" , -- ADDR 1994
			"00000000000000001100110001111001" , -- ADDR 1995
			"00000000000000001010000101111100" , -- ADDR 1996
			"00000000000000001010110101110111" , -- ADDR 1997
			"00000000000000001011011000010111" , -- ADDR 1998
			"00000000000000001000001000010110" , -- ADDR 1999
			"00000000000000001001110101110111" , -- ADDR 2000
			"00000000000000001100000101011001" , -- ADDR 2001
			"00000000000000001001111010100000" , -- ADDR 2002
			"00000000000000010010101101000001" , -- ADDR 2003
			"00000000000000001110000010010001" , -- ADDR 2004
			"00000000000000001000100110011100" , -- ADDR 2005
			"00000000000000001101000000000110" , -- ADDR 2006
			"00000000000000000100110111010101" , -- ADDR 2007
			"00000000000000001101101100010000" , -- ADDR 2008
			"00000000000000001111100000101010" , -- ADDR 2009
			"00000000000000000100101100100011" , -- ADDR 2010
			"00000000000000000101001001100111" , -- ADDR 2011
			"00000000000000001101101010001010" , -- ADDR 2012
			"00000000000000001011111110010001" , -- ADDR 2013
			"00000000000000001100000001100110" , -- ADDR 2014
			"00000000000000010000000011100101" , -- ADDR 2015
			"00000000000000001001010100101000" , -- ADDR 2016
			"00000000000000001011001001010011" , -- ADDR 2017
			"00000000000000001101011110000100" , -- ADDR 2018
			"00000000000000001001010101000010" , -- ADDR 2019
			"00000000000000000110110011110101" , -- ADDR 2020
			"00000000000000001101101111101111" , -- ADDR 2021
			"00000000000000001011000110001101" , -- ADDR 2022
			"00000000000000001110110000011000" , -- ADDR 2023
			"00000000000000001000101000111000" , -- ADDR 2024
			"00000000000000001011110100000000" , -- ADDR 2025
			"00000000000000001010101101010111" , -- ADDR 2026
			"00000000000000001010001010010001" , -- ADDR 2027
			"00000000000000001011101111010011" , -- ADDR 2028
			"00000000000000001110010101000110" , -- ADDR 2029
			"00000000000000001001001011001001" , -- ADDR 2030
			"00000000000000010100011100011010" , -- ADDR 2031
			"00000000000000001111111000011110" , -- ADDR 2032
			"00000000000000001000000001111110" , -- ADDR 2033
			"00000000000000001111000111010111" , -- ADDR 2034
			"00000000000000000101100010010000" , -- ADDR 2035
			"00000000000000001101001001011100" , -- ADDR 2036
			"00000000000000001111000011110101" , -- ADDR 2037
			"00000000000000000100001001101000" , -- ADDR 2038
			"00000000000000001001001101101000" , -- ADDR 2039
			"00000000000000001000010000101110" , -- ADDR 2040
			"00000000000000001101001001011100" , -- ADDR 2041
			"00000000000000001100101000011100" , -- ADDR 2042
			"00000000000000001100101010101100" , -- ADDR 2043
			"00000000000000001010100001100001" , -- ADDR 2044
			"00000000000000001011011110100011" , -- ADDR 2045
			"00000000000000000111110000100100" , -- ADDR 2046
			"00000000000000000111111000110111" , -- ADDR 2047
			"00000000000000001001111000110001" , -- ADDR 2048
			"00000000000000001110101000011101" , -- ADDR 2049
			"00000000000000001100000111110001" , -- ADDR 2050
			"00000000000000001100110011111111" , -- ADDR 2051
			"00000000000000001100000000001011" , -- ADDR 2052
			"00000000000000001101110110010111" , -- ADDR 2053
			"00000000000000000111100010100111" , -- ADDR 2054
			"00000000000000000111000111100011" , -- ADDR 2055
			"00000000000000001001111101100100" , -- ADDR 2056
			"00000000000000001100011011110011" , -- ADDR 2057
			"00000000000000010010011101000111" , -- ADDR 2058
			"00000000000000001101101010001010" , -- ADDR 2059
			"00000000000000001011000100011111" , -- ADDR 2060
			"00000000000000001011111010011011" , -- ADDR 2061
			"00000000000000000011100011100000" , -- ADDR 2062
			"00000000000000010000000100001011" , -- ADDR 2063
			"00000000000000010001110011110001" , -- ADDR 2064
			"00000000000000001001110101110111" , -- ADDR 2065
			"00000000000000000111010100001111" , -- ADDR 2066
			"00000000000000010000011011000100" , -- ADDR 2067
			"00000000000000010000100100111001" , -- ADDR 2068
			"00000000000000001001100010001011" , -- ADDR 2069
			"00000000000000001110011010011010" , -- ADDR 2070
			"00000000000000001111100111101001" , -- ADDR 2071
			"00000000000000001011110100000000" , -- ADDR 2072
			"00000000000000001011000001111001" , -- ADDR 2073
			"00000000000000001101101010100101" , -- ADDR 2074
			"00000000000000001011100011000001" , -- ADDR 2075
			"00000000000000010000010000001101" , -- ADDR 2076
			"00000000000000001101101010100101" , -- ADDR 2077
			"00000000000000001111101001111101" , -- ADDR 2078
			"00000000000000001111110101001110" , -- ADDR 2079
			"00000000000000001011101100001101" , -- ADDR 2080
			"00000000000000001000100110011100" , -- ADDR 2081
			"00000000000000001101001110111011" , -- ADDR 2082
			"00000000000000001110010011100000" , -- ADDR 2083
			"00000000000000010110100110101110" , -- ADDR 2084
			"00000000000000010001110011110001" , -- ADDR 2085
			"00000000000000001101000111010000" , -- ADDR 2086
			"00000000000000001111111100010011" , -- ADDR 2087
			"00000000000000000001000000011011" , -- ADDR 2088
			"00000000000000010010001111101101" , -- ADDR 2089
			"00000000000000010100001000011110" , -- ADDR 2090
			"00000000000000000011101110100000" , -- ADDR 2091
			"00000000000000010100110111000000" , -- ADDR 2092
			"00000000000000001101010010110100" , -- ADDR 2093
			"00000000000000010011000100010110" , -- ADDR 2094
			"00000000000000010000111011101010" , -- ADDR 2095
			"00000000000000001111101101000111" , -- ADDR 2096
			"00000000000000001101110111011110" , -- ADDR 2097
			"00000000000000010000010000101011" , -- ADDR 2098
			"00000000000000001010010001000000" , -- ADDR 2099
			"00000000000000010101000011000001" , -- ADDR 2100
			"00000000000000001110111011001011" , -- ADDR 2101
			"00000000000000010110000001100011" , -- ADDR 2102
			"00000000000000010011000000000011" , -- ADDR 2103
			"00000000000000010110110011111010" , -- ADDR 2104
			"00000000000000001100001100111100" , -- ADDR 2105
			"00000000000000000010100000111000" , -- ADDR 2106
			"00000000000000000111111111110101" , -- ADDR 2107
			"00000000000000010101011110011110" , -- ADDR 2108
			"00000000000000010101010000001100" , -- ADDR 2109
			"00000000000000010000111000111101" , -- ADDR 2110
			"00000000000000010100000100101011" , -- ADDR 2111
			"00000000000000001101011011111100" , -- ADDR 2112
			"00000000000000001000111010010001" , -- ADDR 2113
			"00000000000000011000110111001001" , -- ADDR 2114
			"00000000000000011010011101010110" , -- ADDR 2115
			"00000000000000010101001000001011" , -- ADDR 2116
			"00000000000000001111111001111010" , -- ADDR 2117
			"00000000000000001111111001100011" , -- ADDR 2118
			"00000000000000010001110001001100" , -- ADDR 2119
			"00000000000000010001010101011000" , -- ADDR 2120
			"00000000000000001110101100110000" , -- ADDR 2121
			"00000000000000010000000011100101" , -- ADDR 2122
			"00000000000000001100101111101010" , -- ADDR 2123
			"00000000000000010001110101000011" , -- ADDR 2124
			"00000000000000010000111111010000" , -- ADDR 2125
			"00000000000000010100100110100010" , -- ADDR 2126
			"00000000000000010011100111101010" , -- ADDR 2127
			"00000000000000010110000100111011" , -- ADDR 2128
			"00000000000000001101011101101001" , -- ADDR 2129
			"00000000000000000100100101100100" , -- ADDR 2130
			"00000000000000001010111010110001" , -- ADDR 2131
			"00000000000000010100101000011000" , -- ADDR 2132
			"00000000000000010111100001010010" , -- ADDR 2133
			"00000000000000010010111001100110" , -- ADDR 2134
			"00000000000000010011010010110001" , -- ADDR 2135
			"00000000000000001111110011111001" , -- ADDR 2136
			"00000000000000000110100100101110" , -- ADDR 2137
			"00000000000000011000010100101000" , -- ADDR 2138
			"00000000000000011010000100011100" , -- ADDR 2139
			"00000000000000001101101010100101" , -- ADDR 2140
			"00000000000000010100001000011110" , -- ADDR 2141
			"00000000000000000100101100100011" , -- ADDR 2142
			"00000000000000001000010110011101" , -- ADDR 2143
			"00000000000000000111010000000010" , -- ADDR 2144
			"00000000000000000101011001001011" , -- ADDR 2145
			"00000000000000001101110100011100" , -- ADDR 2146
			"00000000000000010101011001101010" , -- ADDR 2147
			"00000000000000001010100110011001" , -- ADDR 2148
			"00000000000000001001101110010001" , -- ADDR 2149
			"00000000000000000010100011001000" , -- ADDR 2150
			"00000000000000000110000001111010" , -- ADDR 2151
			"00000000000000001001010110010000" , -- ADDR 2152
			"00000000000000010010010110011110" , -- ADDR 2153
			"00000000000000010000001101100000" , -- ADDR 2154
			"00000000000000000110010011001111" , -- ADDR 2155
			"00000000000000001100100000101101" , -- ADDR 2156
			"00000000000000001010000010010110" , -- ADDR 2157
			"00000000000000000101111000010011" , -- ADDR 2158
			"00000000000000001100011011101010" , -- ADDR 2159
			"00000000000000010000010011000001" , -- ADDR 2160
			"00000000000000000110000110111100" , -- ADDR 2161
			"00000000000000000110101101111010" , -- ADDR 2162
			"00000000000000011001000111110111" , -- ADDR 2163
			"00000000000000001001000011110100" , -- ADDR 2164
			"00000000000000000101010110101100" , -- ADDR 2165
			"00000000000000000111110110001100" , -- ADDR 2166
			"00000000000000001100011111010101" , -- ADDR 2167
			"00000000000000000011001011001000" , -- ADDR 2168
			"00000000000000011011000001010011" , -- ADDR 2169
			"00000000000000000011001011101110" , -- ADDR 2170
			"00000000000000010100100101000011" , -- ADDR 2171
			"00000000000000001011000111100101" , -- ADDR 2172
			"00000000000000010010101011110011" , -- ADDR 2173
			"00000000000000000110000110101000" , -- ADDR 2174
			"00000000000000001011010111101101" , -- ADDR 2175
			"00000000000000000101010111110000" , -- ADDR 2176
			"00000000000000010010000101001101" , -- ADDR 2177
			"00000000000000001000000111011010" , -- ADDR 2178
			"00000000000000000100101100001001" , -- ADDR 2179
			"00000000000000010000110110001000" , -- ADDR 2180
			"00000000000000000001001111101011" , -- ADDR 2181
			"00000000000000001111101110111100" , -- ADDR 2182
			"00000000000000010011100110011001" , -- ADDR 2183
			"00000000000000010100011000011111" , -- ADDR 2184
			"00000000000000010100010000111110" , -- ADDR 2185
			"00000000000000010110110010100101" , -- ADDR 2186
			"00000000000000010010101001011101" , -- ADDR 2187
			"00000000000000001111100101000100" , -- ADDR 2188
			"00000000000000010110100001111010" , -- ADDR 2189
			"00000000000000000010000000110110" , -- ADDR 2190
			"00000000000000011000000010111110" , -- ADDR 2191
			"00000000000000001100011101000010" , -- ADDR 2192
			"00000000000000010100100011111100" , -- ADDR 2193
			"00000000000000010000100000010010" , -- ADDR 2194
			"00000000000000010011011010010111" , -- ADDR 2195
			"00000000000000010010000110100100" , -- ADDR 2196
			"00000000000000010110100010010101" , -- ADDR 2197
			"00000000000000001111001000100000" , -- ADDR 2198
			"00000000000000011101101111100100" , -- ADDR 2199
			"00000000000000011001001101000110" , -- ADDR 2200
			"00000000000000001110101100000110" , -- ADDR 2201
			"00000000000000011000010001001011" , -- ADDR 2202
			"00000000000000001010100010100110" , -- ADDR 2203
			"00000000000000010010111000000110" , -- ADDR 2204
			"00000000000000010100110011011100" , -- ADDR 2205
			"00000000000000000011111010000000" , -- ADDR 2206
			"00000000000000000011000101101001" , -- ADDR 2207
			"00000000000000000100110110001001" , -- ADDR 2208
			"00000000000000001001001001000011" , -- ADDR 2209
			"00000000000000010101110110011011" , -- ADDR 2210
			"00000000000000000110000111111000" , -- ADDR 2211
			"00000000000000001100010110100100" , -- ADDR 2212
			"00000000000000000010010000000100" , -- ADDR 2213
			"00000000000000001001110001000000" , -- ADDR 2214
			"00000000000000000100111000100000" , -- ADDR 2215
			"00000000000000001110011011010101" , -- ADDR 2216
			"00000000000000001011100110010100" , -- ADDR 2217
			"00000000000000001001011001000111" , -- ADDR 2218
			"00000000000000001001110001000000" , -- ADDR 2219
			"00000000000000000110000010100011" , -- ADDR 2220
			"00000000000000001000010110011101" , -- ADDR 2221
			"00000000000000000111110100010000" , -- ADDR 2222
			"00000000000000001110000001010100" , -- ADDR 2223
			"00000000000000001010100010100110" , -- ADDR 2224
			"00000000000000001011011000010111" , -- ADDR 2225
			"00000000000000000100001001001011" , -- ADDR 2226
			"00000000000000001000001101001111" , -- ADDR 2227
			"00000000000000000110010011001111" , -- ADDR 2228
			"00000000000000011000100001100001" , -- ADDR 2229
			"00000000000000000010010000000100" , -- ADDR 2230
			"00000000000000010000000110110010" , -- ADDR 2231
			"00000000000000000101110011011010" , -- ADDR 2232
			"00000000000000001101101011000000" , -- ADDR 2233
			"00000000000000000100000001101100" , -- ADDR 2234
			"00000000000000001101010100111101" , -- ADDR 2235
			"00000000000000001001000000011100" , -- ADDR 2236
			"00000000000000001101010000111100" , -- ADDR 2237
			"00000000000000000111000010101100" , -- ADDR 2238
			"00000000000000000010011100010000" , -- ADDR 2239
			"00000000000000001100001010011100" , -- ADDR 2240
			"00000000000000000100001001101000" , -- ADDR 2241
			"00000000000000001111000000011001" , -- ADDR 2242
			"00000000000000001110010111101000" , -- ADDR 2243
			"00000000000000001111000011110101" , -- ADDR 2244
			"00000000000000000100101001010010" , -- ADDR 2245
			"00000000000000000110111100101100" , -- ADDR 2246
			"00000000000000010100011000011111" , -- ADDR 2247
			"00000000000000000101101011011011" , -- ADDR 2248
			"00000000000000001100101110111010" , -- ADDR 2249
			"00000000000000000101001001100111" , -- ADDR 2250
			"00000000000000001011001000100111" , -- ADDR 2251
			"00000000000000000010001011110000" , -- ADDR 2252
			"00000000000000001011010110110111" , -- ADDR 2253
			"00000000000000001001000101100000" , -- ADDR 2254
			"00000000000000001010010110111010" , -- ADDR 2255
			"00000000000000001011001000100111" , -- ADDR 2256
			"00000000000000000110100100011011" , -- ADDR 2257
			"00000000000000001001000100000001" , -- ADDR 2258
			"00000000000000000110101010011111" , -- ADDR 2259
			"00000000000000001011010011110101" , -- ADDR 2260
			"00000000000000001100011100101110" , -- ADDR 2261
			"00000000000000001101100111001110" , -- ADDR 2262
			"00000000000000001011011001100010" , -- ADDR 2263
			"00000000000000010001000101110000" , -- ADDR 2264
			"00000000000000001010001000001101" , -- ADDR 2265
			"00000000000000001000000101110000" , -- ADDR 2266
			"00000000000000000101000010001000" , -- ADDR 2267
			"00000000000000000110111000010010" , -- ADDR 2268
			"00000000000000000110101000011110" , -- ADDR 2269
			"00000000000000001101110100001010" , -- ADDR 2270
			"00000000000000001101001101000011" , -- ADDR 2271
			"00000000000000000101110111101010" , -- ADDR 2272
			"00000000000000001110100110101000" , -- ADDR 2273
			"00000000000000001010100101110110" , -- ADDR 2274
			"00000000000000000100100000000111" , -- ADDR 2275
			"00000000000000001011010010111111" , -- ADDR 2276
			"00000000000000001010111010110001" , -- ADDR 2277
			"00000000000000001000101010001100" , -- ADDR 2278
			"00000000000000001010001100101101" , -- ADDR 2279
			"00000000000000011000011110010000" , -- ADDR 2280
			"00000000000000000100110111010101" , -- ADDR 2281
			"00000000000000010011010100110110" , -- ADDR 2282
			"00000000000000001011011000010111" , -- ADDR 2283
			"00000000000000010010000100111001" , -- ADDR 2284
			"00000000000000000100110010111111" , -- ADDR 2285
			"00000000000000001000001111000110" , -- ADDR 2286
			"00000000000000000010101110101100" , -- ADDR 2287
			"00000000000000010001001111010100" , -- ADDR 2288
			"00000000000000001010111111010011" , -- ADDR 2289
			"00000000000000000110110011110101" , -- ADDR 2290
			"00000000000000001111111001011011" , -- ADDR 2291
			"00000000000000000011001011001000" , -- ADDR 2292
			"00000000000000001100110001111001" , -- ADDR 2293
			"00000000000000010011010111001110" , -- ADDR 2294
			"00000000000000010100011011000000" , -- ADDR 2295
			"00000000000000011001110110100011" , -- ADDR 2296
			"00000000000000001101000111111111" , -- ADDR 2297
			"00000000000000010110000000011011" , -- ADDR 2298
			"00000000000000010001010110010111" , -- ADDR 2299
			"00000000000000010101001111011110" , -- ADDR 2300
			"00000000000000010100000111001001" , -- ADDR 2301
			"00000000000000011000100001110000" , -- ADDR 2302
			"00000000000000010000000100001011" , -- ADDR 2303
			"00000000000000011111011011010101" , -- ADDR 2304
			"00000000000000011010111100110110" , -- ADDR 2305
			"00000000000000001111110001101110" , -- ADDR 2306
			"00000000000000011010001001000011" , -- ADDR 2307
			"00000000000000001100100011011100" , -- ADDR 2308
			"00000000000000010011101000011011" , -- ADDR 2309
			"00000000000000010101100000110111" , -- ADDR 2310
			"00000000000000010010001001011010" , -- ADDR 2311
			"00000000000000001000000011011001" , -- ADDR 2312
			"00000000000000001111111000000111" , -- ADDR 2313
			"00000000000000000100101010100001" , -- ADDR 2314
			"00000000000000001100101100101010" , -- ADDR 2315
			"00000000000000000111100100101000" , -- ADDR 2316
			"00000000000000001111011010010111" , -- ADDR 2317
			"00000000000000000110100100101110" , -- ADDR 2318
			"00000000000000000001111101111110" , -- ADDR 2319
			"00000000000000001110010000110101" , -- ADDR 2320
			"00000000000000000010000100100101" , -- ADDR 2321
			"00000000000000001111100010010000" , -- ADDR 2322
			"00000000000000010000100111100010" , -- ADDR 2323
			"00000000000000010001010011100000" , -- ADDR 2324
			"00000000000000001011010111000010" , -- ADDR 2325
			"00000000000000000100010111100001" , -- ADDR 2326
			"00000000000000001110101001100000" , -- ADDR 2327
			"00000000000000010011111000000101" , -- ADDR 2328
			"00000000000000010100110101010001" , -- ADDR 2329
			"00000000000000000011011100111110" , -- ADDR 2330
			"00000000000000010101110101100011" , -- ADDR 2331
			"00000000000000010010011000010110" , -- ADDR 2332
			"00000000000000000100000010101001" , -- ADDR 2333
			"00000000000000010011011000101100" , -- ADDR 2334
			"00000000000000001110001001111111" , -- ADDR 2335
			"00000000000000000110100000111011" , -- ADDR 2336
			"00000000000000001000011000111110" , -- ADDR 2337
			"00000000000000001000001100000101" , -- ADDR 2338
			"00000000000000000111000110001101" , -- ADDR 2339
			"00000000000000010000011111001111" , -- ADDR 2340
			"00000000000000001101110110010111" , -- ADDR 2341
			"00000000000000001000000111011010" , -- ADDR 2342
			"00000000000000001010011111001001" , -- ADDR 2343
			"00000000000000000111100100011000" , -- ADDR 2344
			"00000000000000000111010101000001" , -- ADDR 2345
			"00000000000000001001111000110001" , -- ADDR 2346
			"00000000000000001111011000011000" , -- ADDR 2347
			"00000000000000001000100110011100" , -- ADDR 2348
			"00000000000000001001010000111011" , -- ADDR 2349
			"00000000000000001101010010000110" , -- ADDR 2350
			"00000000000000010100011100011010" , -- ADDR 2351
			"00000000000000010100000010011111" , -- ADDR 2352
			"00000000000000000001100010110101" , -- ADDR 2353
			"00000000000000010010100001110111" , -- ADDR 2354
			"00000000000000001111101100011001" , -- ADDR 2355
			"00000000000000000010110010001010" , -- ADDR 2356
			"00000000000000010001011100011001" , -- ADDR 2357
			"00000000000000010000000101000111" , -- ADDR 2358
			"00000000000000000010011111010110" , -- ADDR 2359
			"00000000000000000100011101001000" , -- ADDR 2360
			"00000000000000001001101110101010" , -- ADDR 2361
			"00000000000000000110111010001110" , -- ADDR 2362
			"00000000000000001100011100101110" , -- ADDR 2363
			"00000000000000001010111010110001" , -- ADDR 2364
			"00000000000000000110000111100100" , -- ADDR 2365
			"00000000000000001011000111100101" , -- ADDR 2366
			"00000000000000000101000010001000" , -- ADDR 2367
			"00000000000000001011000010000100" , -- ADDR 2368
			"00000000000000001110101000011101" , -- ADDR 2369
			"00000000000000001111110010010101" , -- ADDR 2370
			"00000000000000000110010101010110" , -- ADDR 2371
			"00000000000000010011001001001001" , -- ADDR 2372
			"00000000000000010011001001001001" , -- ADDR 2373
			"00000000000000001110101001100000" , -- ADDR 2374
			"00000000000000010001101110101110" , -- ADDR 2375
			"00000000000000001011010111000010" , -- ADDR 2376
			"00000000000000000111100110101001" , -- ADDR 2377
			"00000000000000010110011100011111" , -- ADDR 2378
			"00000000000000011000000000101111" , -- ADDR 2379
			"00000000000000010011000100011101" , -- ADDR 2380
			"00000000000000001101011101101001" , -- ADDR 2381
			"00000000000000001001011111110001" , -- ADDR 2382
			"00000000000000010001101011100110" , -- ADDR 2383
			"00000000000000000101101111110001" , -- ADDR 2384
			"00000000000000001100010001001001" , -- ADDR 2385
			"00000000000000010101100000110111" , -- ADDR 2386
			"00000000000000010110101100100010" , -- ADDR 2387
			"00000000000000010010100101111110" , -- ADDR 2388
			"00000000000000001111011010101111" , -- ADDR 2389
			"00000000000000000001011011000111" , -- ADDR 2390
			"00000000000000010000110110100101" , -- ADDR 2391
			"00000000000000001110100100100010" , -- ADDR 2392
			"00000000000000000100000001101100" , -- ADDR 2393
			"00000000000000000101111111000011" , -- ADDR 2394
			"00000000000000000100110011110010" , -- ADDR 2395
			"00000000000000010001110011000001" , -- ADDR 2396
			"00000000000000000111110100010000" , -- ADDR 2397
			"00000000000000010101111100101100" , -- ADDR 2398
			"00000000000000010010011000110001" , -- ADDR 2399
			"00000000000000010010010111101000" , -- ADDR 2400
			"00000000000000001110011000111101" , -- ADDR 2401
			"00000000000000000011110100100100" , -- ADDR 2402
			"00000000000000010001001001000110" , -- ADDR 2403
			"00000000000000010000001001001001" , -- ADDR 2404
			"00000000000000010000100111100010" , -- ADDR 2405
			"00000000000000001111101000001000" , -- ADDR 2406
			"00000000000000001101010100111101" , -- ADDR 2407
			"00000000000000000101001000100000" , -- ADDR 2408
			"00000000000000000111000001111000" , -- ADDR 2409
			"00000000000000001111001000111000" , -- ADDR 2410
			"00000000000000010010010110110010" , -- ADDR 2411
			"00000000000000010011001001100011" , -- ADDR 2412
			"00000000000000010010011101000111" , -- ADDR 2413
			"00000000000000010100010011111001" , -- ADDR 2414
			"00000000000000000001111101111110" , -- ADDR 2415
			"00000000000000000000000000000000" , -- ADDR 2416
			"00000000000000000000000000000000" , -- ADDR 2417
			"00000000000000000000000000000000" , -- ADDR 2418
			"00000000000000000000000000000000" , -- ADDR 2419
			"00000000000000000000000000000000" , -- ADDR 2420
			"00000000000000000000000000000000" , -- ADDR 2421
			"00000000000000000000000000000000" , -- ADDR 2422
			"00000000000000000000000000000000" , -- ADDR 2423
			"00000000000000000000000000000000" , -- ADDR 2424
			"00000000000000000000000000000000" , -- ADDR 2425
			"00000000000000000000000000000000" , -- ADDR 2426
			"00000000000000000000000000000000" , -- ADDR 2427
			"00000000000000000000000000000000" , -- ADDR 2428
			"00000000000000000000000000000000" , -- ADDR 2429
			"00000000000000000000000000000000" , -- ADDR 2430
			"00000000000000000000000000000000" , -- ADDR 2431
			"00000000000000000000000000000000" , -- ADDR 2432
			"00000000000000000000000000000000" , -- ADDR 2433
			"00000000000000000000000000000000" , -- ADDR 2434
			"00000000000000000000000000000000" , -- ADDR 2435
			"00000000000000000000000000000000" , -- ADDR 2436
			"00000000000000000000000000000000" , -- ADDR 2437
			"00000000000000000000000000000000" , -- ADDR 2438
			"00000000000000000000000000000000" , -- ADDR 2439
			"00000000000000000000000000000000" , -- ADDR 2440
			"00000000000000000000000000000000" , -- ADDR 2441
			"00000000000000000000000000000000" , -- ADDR 2442
			"00000000000000000000000000000000" , -- ADDR 2443
			"00000000000000000000000000000000" , -- ADDR 2444
			"00000000000000000000000000000000" , -- ADDR 2445
			"00000000000000000000000000000000" , -- ADDR 2446
			"00000000000000000000000000000000" , -- ADDR 2447
			"00000000000000000000000000000000" , -- ADDR 2448
			"00000000000000000000000000000000" , -- ADDR 2449
			"00000000000000000000000000000000" , -- ADDR 2450
			"00000000000000000000000000000000" , -- ADDR 2451
			"00000000000000000000000000000000" , -- ADDR 2452
			"00000000000000000000000000000000" , -- ADDR 2453
			"00000000000000000000000000000000" , -- ADDR 2454
			"00000000000000000000000000000000" , -- ADDR 2455
			"00000000000000000000000000000000" , -- ADDR 2456
			"00000000000000000000000000000000" , -- ADDR 2457
			"00000000000000000000000000000000" , -- ADDR 2458
			"00000000000000000000000000000000" , -- ADDR 2459
			"00000000000000000000000000000000" , -- ADDR 2460
			"00000000000000000000000000000000" , -- ADDR 2461
			"00000000000000000000000000000000" , -- ADDR 2462
			"00000000000000000000000000000000" , -- ADDR 2463
			"00000000000000000000000000000000" , -- ADDR 2464
			"00000000000000000000000000000000" , -- ADDR 2465
			"00000000000000000000000000000000" , -- ADDR 2466
			"00000000000000000000000000000000" , -- ADDR 2467
			"00000000000000000000000000000000" , -- ADDR 2468
			"00000000000000000000000000000000" , -- ADDR 2469
			"00000000000000000000000000000000" , -- ADDR 2470
			"00000000000000000000000000000000" , -- ADDR 2471
			"00000000000000000000000000000000" , -- ADDR 2472
			"00000000000000000000000000000000" , -- ADDR 2473
			"00000000000000000000000000000000" , -- ADDR 2474
			"00000000000000000000000000000000" , -- ADDR 2475
			"00000000000000000000000000000000" , -- ADDR 2476
			"00000000000000000000000000000000" , -- ADDR 2477
			"00000000000000000000000000000000" , -- ADDR 2478
			"00000000000000000000000000000000" , -- ADDR 2479
			"00000000000000000000000000000000" , -- ADDR 2480
			"00000000000000000000000000000000" , -- ADDR 2481
			"00000000000000000000000000000000" , -- ADDR 2482
			"00000000000000000000000000000000" , -- ADDR 2483
			"00000000000000000000000000000000" , -- ADDR 2484
			"00000000000000000000000000000000" , -- ADDR 2485
			"00000000000000000000000000000000" , -- ADDR 2486
			"00000000000000000000000000000000" , -- ADDR 2487
			"00000000000000000000000000000000" , -- ADDR 2488
			"00000000000000000000000000000000" , -- ADDR 2489
			"00000000000000000000000000000000" , -- ADDR 2490
			"00000000000000000000000000000000" , -- ADDR 2491
			"00000000000000000000000000000000" , -- ADDR 2492
			"00000000000000000000000000000000" , -- ADDR 2493
			"00000000000000000000000000000000" , -- ADDR 2494
			"00000000000000000000000000000000" , -- ADDR 2495
			"00000000000000000000000000000000" , -- ADDR 2496
			"00000000000000000000000000000000" , -- ADDR 2497
			"00000000000000000000000000000000" , -- ADDR 2498
			"00000000000000000000000000000000" , -- ADDR 2499
			"00000000000000000000000000000000" , -- ADDR 2500
			"00000000000000000000000000000000" , -- ADDR 2501
			"00000000000000000000000000000000" , -- ADDR 2502
			"00000000000000000000000000000000" , -- ADDR 2503
			"00000000000000000000000000000000" , -- ADDR 2504
			"00000000000000000000000000000000" , -- ADDR 2505
			"00000000000000000000000000000000" , -- ADDR 2506
			"00000000000000000000000000000000" , -- ADDR 2507
			"00000000000000000000000000000000" , -- ADDR 2508
			"00000000000000000000000000000000" , -- ADDR 2509
			"00000000000000000000000000000000" , -- ADDR 2510
			"00000000000000000000000000000000" , -- ADDR 2511
			"00000000000000000000000000000000" , -- ADDR 2512
			"00000000000000000000000000000000" , -- ADDR 2513
			"00000000000000000000000000000000" , -- ADDR 2514
			"00000000000000000000000000000000" , -- ADDR 2515
			"00000000000000000000000000000000" , -- ADDR 2516
			"00000000000000000000000000000000" , -- ADDR 2517
			"00000000000000000000000000000000" , -- ADDR 2518
			"00000000000000000000000000000000" , -- ADDR 2519
			"00000000000000000000000000000000" , -- ADDR 2520
			"00000000000000000000000000000000" , -- ADDR 2521
			"00000000000000000000000000000000" , -- ADDR 2522
			"00000000000000000000000000000000" , -- ADDR 2523
			"00000000000000000000000000000000" , -- ADDR 2524
			"00000000000000000000000000000000" , -- ADDR 2525
			"00000000000000000000000000000000" , -- ADDR 2526
			"00000000000000000000000000000000" , -- ADDR 2527
			"00000000000000000000000000000000" , -- ADDR 2528
			"00000000000000000000000000000000" , -- ADDR 2529
			"00000000000000000000000000000000" , -- ADDR 2530
			"00000000000000000000000000000000" , -- ADDR 2531
			"00000000000000000000000000000000" , -- ADDR 2532
			"00000000000000000000000000000000" , -- ADDR 2533
			"00000000000000000000000000000000" , -- ADDR 2534
			"00000000000000000000000000000000" , -- ADDR 2535
			"00000000000000000000000000000000" , -- ADDR 2536
			"00000000000000000000000000000000" , -- ADDR 2537
			"00000000000000000000000000000000" , -- ADDR 2538
			"00000000000000000000000000000000" , -- ADDR 2539
			"00000000000000000000000000000000" , -- ADDR 2540
			"00000000000000000000000000000000" , -- ADDR 2541
			"00000000000000000000000000000000" , -- ADDR 2542
			"00000000000000000000000000000000" , -- ADDR 2543
			"00000000000000000000000000000000" , -- ADDR 2544
			"00000000000000000000000000000000" , -- ADDR 2545
			"00000000000000000000000000000000" , -- ADDR 2546
			"00000000000000000000000000000000" , -- ADDR 2547
			"00000000000000000000000000000000" , -- ADDR 2548
			"00000000000000000000000000000000" , -- ADDR 2549
			"00000000000000000000000000000000" , -- ADDR 2550
			"00000000000000000000000000000000" , -- ADDR 2551
			"00000000000000000000000000000000" , -- ADDR 2552
			"00000000000000000000000000000000" , -- ADDR 2553
			"00000000000000000000000000000000" , -- ADDR 2554
			"00000000000000000000000000000000" , -- ADDR 2555
			"00000000000000000000000000000000" , -- ADDR 2556
			"00000000000000000000000000000000" , -- ADDR 2557
			"00000000000000000000000000000000" , -- ADDR 2558
			"00000000000000000000000000000000" , -- ADDR 2559
			"00000000000000000000000000000000" , -- ADDR 2560
			"00000000000000000000000000000000" , -- ADDR 2561
			"00000000000000000000000000000000" , -- ADDR 2562
			"00000000000000000000000000000000" , -- ADDR 2563
			"00000000000000000000000000000000" , -- ADDR 2564
			"00000000000000000000000000000000" , -- ADDR 2565
			"00000000000000000000000000000000" , -- ADDR 2566
			"00000000000000000000000000000000" , -- ADDR 2567
			"00000000000000000000000000000000" , -- ADDR 2568
			"00000000000000000000000000000000" , -- ADDR 2569
			"00000000000000000000000000000000" , -- ADDR 2570
			"00000000000000000000000000000000" , -- ADDR 2571
			"00000000000000000000000000000000" , -- ADDR 2572
			"00000000000000000000000000000000" , -- ADDR 2573
			"00000000000000000000000000000000" , -- ADDR 2574
			"00000000000000000000000000000000" , -- ADDR 2575
			"00000000000000000000000000000000" , -- ADDR 2576
			"00000000000000000000000000000000" , -- ADDR 2577
			"00000000000000000000000000000000" , -- ADDR 2578
			"00000000000000000000000000000000" , -- ADDR 2579
			"00000000000000000000000000000000" , -- ADDR 2580
			"00000000000000000000000000000000" , -- ADDR 2581
			"00000000000000000000000000000000" , -- ADDR 2582
			"00000000000000000000000000000000" , -- ADDR 2583
			"00000000000000000000000000000000" , -- ADDR 2584
			"00000000000000000000000000000000" , -- ADDR 2585
			"00000000000000000000000000000000" , -- ADDR 2586
			"00000000000000000000000000000000" , -- ADDR 2587
			"00000000000000000000000000000000" , -- ADDR 2588
			"00000000000000000000000000000000" , -- ADDR 2589
			"00000000000000000000000000000000" , -- ADDR 2590
			"00000000000000000000000000000000" , -- ADDR 2591
			"00000000000000000000000000000000" , -- ADDR 2592
			"00000000000000000000000000000000" , -- ADDR 2593
			"00000000000000000000000000000000" , -- ADDR 2594
			"00000000000000000000000000000000" , -- ADDR 2595
			"00000000000000000000000000000000" , -- ADDR 2596
			"00000000000000000000000000000000" , -- ADDR 2597
			"00000000000000000000000000000000" , -- ADDR 2598
			"00000000000000000000000000000000" , -- ADDR 2599
			"00000000000000000000000000000000" , -- ADDR 2600
			"00000000000000000000000000000000" , -- ADDR 2601
			"00000000000000000000000000000000" , -- ADDR 2602
			"00000000000000000000000000000000" , -- ADDR 2603
			"00000000000000000000000000000000" , -- ADDR 2604
			"00000000000000000000000000000000" , -- ADDR 2605
			"00000000000000000000000000000000" , -- ADDR 2606
			"00000000000000000000000000000000" , -- ADDR 2607
			"00000000000000000000000000000000" , -- ADDR 2608
			"00000000000000000000000000000000" , -- ADDR 2609
			"00000000000000000000000000000000" , -- ADDR 2610
			"00000000000000000000000000000000" , -- ADDR 2611
			"00000000000000000000000000000000" , -- ADDR 2612
			"00000000000000000000000000000000" , -- ADDR 2613
			"00000000000000000000000000000000" , -- ADDR 2614
			"00000000000000000000000000000000" , -- ADDR 2615
			"00000000000000000000000000000000" , -- ADDR 2616
			"00000000000000000000000000000000" , -- ADDR 2617
			"00000000000000000000000000000000" , -- ADDR 2618
			"00000000000000000000000000000000" , -- ADDR 2619
			"00000000000000000000000000000000" , -- ADDR 2620
			"00000000000000000000000000000000" , -- ADDR 2621
			"00000000000000000000000000000000" , -- ADDR 2622
			"00000000000000000000000000000000" , -- ADDR 2623
			"00000000000000000000000000000000" , -- ADDR 2624
			"00000000000000000000000000000000" , -- ADDR 2625
			"00000000000000000000000000000000" , -- ADDR 2626
			"00000000000000000000000000000000" , -- ADDR 2627
			"00000000000000000000000000000000" , -- ADDR 2628
			"00000000000000000000000000000000" , -- ADDR 2629
			"00000000000000000000000000000000" , -- ADDR 2630
			"00000000000000000000000000000000" , -- ADDR 2631
			"00000000000000000000000000000000" , -- ADDR 2632
			"00000000000000000000000000000000" , -- ADDR 2633
			"00000000000000000000000000000000" , -- ADDR 2634
			"00000000000000000000000000000000" , -- ADDR 2635
			"00000000000000000000000000000000" , -- ADDR 2636
			"00000000000000000000000000000000" , -- ADDR 2637
			"00000000000000000000000000000000" , -- ADDR 2638
			"00000000000000000000000000000000" , -- ADDR 2639
			"00000000000000000000000000000000" , -- ADDR 2640
			"00000000000000000000000000000000" , -- ADDR 2641
			"00000000000000000000000000000000" , -- ADDR 2642
			"00000000000000000000000000000000" , -- ADDR 2643
			"00000000000000000000000000000000" , -- ADDR 2644
			"00000000000000000000000000000000" , -- ADDR 2645
			"00000000000000000000000000000000" , -- ADDR 2646
			"00000000000000000000000000000000" , -- ADDR 2647
			"00000000000000000000000000000000" , -- ADDR 2648
			"00000000000000000000000000000000" , -- ADDR 2649
			"00000000000000000000000000000000" , -- ADDR 2650
			"00000000000000000000000000000000" , -- ADDR 2651
			"00000000000000000000000000000000" , -- ADDR 2652
			"00000000000000000000000000000000" , -- ADDR 2653
			"00000000000000000000000000000000" , -- ADDR 2654
			"00000000000000000000000000000000" , -- ADDR 2655
			"00000000000000000000000000000000" , -- ADDR 2656
			"00000000000000000000000000000000" , -- ADDR 2657
			"00000000000000000000000000000000" , -- ADDR 2658
			"00000000000000000000000000000000" , -- ADDR 2659
			"00000000000000000000000000000000" , -- ADDR 2660
			"00000000000000000000000000000000" , -- ADDR 2661
			"00000000000000000000000000000000" , -- ADDR 2662
			"00000000000000000000000000000000" , -- ADDR 2663
			"00000000000000000000000000000000" , -- ADDR 2664
			"00000000000000000000000000000000" , -- ADDR 2665
			"00000000000000000000000000000000" , -- ADDR 2666
			"00000000000000000000000000000000" , -- ADDR 2667
			"00000000000000000000000000000000" , -- ADDR 2668
			"00000000000000000000000000000000" , -- ADDR 2669
			"00000000000000000000000000000000" , -- ADDR 2670
			"00000000000000000000000000000000" , -- ADDR 2671
			"00000000000000000000000000000000" , -- ADDR 2672
			"00000000000000000000000000000000" , -- ADDR 2673
			"00000000000000000000000000000000" , -- ADDR 2674
			"00000000000000000000000000000000" , -- ADDR 2675
			"00000000000000000000000000000000" , -- ADDR 2676
			"00000000000000000000000000000000" , -- ADDR 2677
			"00000000000000000000000000000000" , -- ADDR 2678
			"00000000000000000000000000000000" , -- ADDR 2679
			"00000000000000000000000000000000" , -- ADDR 2680
			"00000000000000000000000000000000" , -- ADDR 2681
			"00000000000000000000000000000000" , -- ADDR 2682
			"00000000000000000000000000000000" , -- ADDR 2683
			"00000000000000000000000000000000" , -- ADDR 2684
			"00000000000000000000000000000000" , -- ADDR 2685
			"00000000000000000000000000000000" , -- ADDR 2686
			"00000000000000000000000000000000" , -- ADDR 2687
			"00000000000000000000000000000000" , -- ADDR 2688
			"00000000000000000000000000000000" , -- ADDR 2689
			"00000000000000000000000000000000" , -- ADDR 2690
			"00000000000000000000000000000000" , -- ADDR 2691
			"00000000000000000000000000000000" , -- ADDR 2692
			"00000000000000000000000000000000" , -- ADDR 2693
			"00000000000000000000000000000000" , -- ADDR 2694
			"00000000000000000000000000000000" , -- ADDR 2695
			"00000000000000000000000000000000" , -- ADDR 2696
			"00000000000000000000000000000000" , -- ADDR 2697
			"00000000000000000000000000000000" , -- ADDR 2698
			"00000000000000000000000000000000" , -- ADDR 2699
			"00000000000000000000000000000000" , -- ADDR 2700
			"00000000000000000000000000000000" , -- ADDR 2701
			"00000000000000000000000000000000" , -- ADDR 2702
			"00000000000000000000000000000000" , -- ADDR 2703
			"00000000000000000000000000000000" , -- ADDR 2704
			"00000000000000000000000000000000" , -- ADDR 2705
			"00000000000000000000000000000000" , -- ADDR 2706
			"00000000000000000000000000000000" , -- ADDR 2707
			"00000000000000000000000000000000" , -- ADDR 2708
			"00000000000000000000000000000000" , -- ADDR 2709
			"00000000000000000000000000000000" , -- ADDR 2710
			"00000000000000000000000000000000" , -- ADDR 2711
			"00000000000000000000000000000000" , -- ADDR 2712
			"00000000000000000000000000000000" , -- ADDR 2713
			"00000000000000000000000000000000" , -- ADDR 2714
			"00000000000000000000000000000000" , -- ADDR 2715
			"00000000000000000000000000000000" , -- ADDR 2716
			"00000000000000000000000000000000" , -- ADDR 2717
			"00000000000000000000000000000000" , -- ADDR 2718
			"00000000000000000000000000000000" , -- ADDR 2719
			"00000000000000000000000000000000" , -- ADDR 2720
			"00000000000000000000000000000000" , -- ADDR 2721
			"00000000000000000000000000000000" , -- ADDR 2722
			"00000000000000000000000000000000" , -- ADDR 2723
			"00000000000000000000000000000000" , -- ADDR 2724
			"00000000000000000000000000000000" , -- ADDR 2725
			"00000000000000000000000000000000" , -- ADDR 2726
			"00000000000000000000000000000000" , -- ADDR 2727
			"00000000000000000000000000000000" , -- ADDR 2728
			"00000000000000000000000000000000" , -- ADDR 2729
			"00000000000000000000000000000000" , -- ADDR 2730
			"00000000000000000000000000000000" , -- ADDR 2731
			"00000000000000000000000000000000" , -- ADDR 2732
			"00000000000000000000000000000000" , -- ADDR 2733
			"00000000000000000000000000000000" , -- ADDR 2734
			"00000000000000000000000000000000" , -- ADDR 2735
			"00000000000000000000000000000000" , -- ADDR 2736
			"00000000000000000000000000000000" , -- ADDR 2737
			"00000000000000000000000000000000" , -- ADDR 2738
			"00000000000000000000000000000000" , -- ADDR 2739
			"00000000000000000000000000000000" , -- ADDR 2740
			"00000000000000000000000000000000" , -- ADDR 2741
			"00000000000000000000000000000000" , -- ADDR 2742
			"00000000000000000000000000000000" , -- ADDR 2743
			"00000000000000000000000000000000" , -- ADDR 2744
			"00000000000000000000000000000000" , -- ADDR 2745
			"00000000000000000000000000000000" , -- ADDR 2746
			"00000000000000000000000000000000" , -- ADDR 2747
			"00000000000000000000000000000000" , -- ADDR 2748
			"00000000000000000000000000000000" , -- ADDR 2749
			"00000000000000000000000000000000" , -- ADDR 2750
			"00000000000000000000000000000000" , -- ADDR 2751
			"00000000000000000000000000000000" , -- ADDR 2752
			"00000000000000000000000000000000" , -- ADDR 2753
			"00000000000000000000000000000000" , -- ADDR 2754
			"00000000000000000000000000000000" , -- ADDR 2755
			"00000000000000000000000000000000" , -- ADDR 2756
			"00000000000000000000000000000000" , -- ADDR 2757
			"00000000000000000000000000000000" , -- ADDR 2758
			"00000000000000000000000000000000" , -- ADDR 2759
			"00000000000000000000000000000000" , -- ADDR 2760
			"00000000000000000000000000000000" , -- ADDR 2761
			"00000000000000000000000000000000" , -- ADDR 2762
			"00000000000000000000000000000000" , -- ADDR 2763
			"00000000000000000000000000000000" , -- ADDR 2764
			"00000000000000000000000000000000" , -- ADDR 2765
			"00000000000000000000000000000000" , -- ADDR 2766
			"00000000000000000000000000000000" , -- ADDR 2767
			"00000000000000000000000000000000" , -- ADDR 2768
			"00000000000000000000000000000000" , -- ADDR 2769
			"00000000000000000000000000000000" , -- ADDR 2770
			"00000000000000000000000000000000" , -- ADDR 2771
			"00000000000000000000000000000000" , -- ADDR 2772
			"00000000000000000000000000000000" , -- ADDR 2773
			"00000000000000000000000000000000" , -- ADDR 2774
			"00000000000000000000000000000000" , -- ADDR 2775
			"00000000000000000000000000000000" , -- ADDR 2776
			"00000000000000000000000000000000" , -- ADDR 2777
			"00000000000000000000000000000000" , -- ADDR 2778
			"00000000000000000000000000000000" , -- ADDR 2779
			"00000000000000000000000000000000" , -- ADDR 2780
			"00000000000000000000000000000000" , -- ADDR 2781
			"00000000000000000000000000000000" , -- ADDR 2782
			"00000000000000000000000000000000" , -- ADDR 2783
			"00000000000000000000000000000000" , -- ADDR 2784
			"00000000000000000000000000000000" , -- ADDR 2785
			"00000000000000000000000000000000" , -- ADDR 2786
			"00000000000000000000000000000000" , -- ADDR 2787
			"00000000000000000000000000000000" , -- ADDR 2788
			"00000000000000000000000000000000" , -- ADDR 2789
			"00000000000000000000000000000000" , -- ADDR 2790
			"00000000000000000000000000000000" , -- ADDR 2791
			"00000000000000000000000000000000" , -- ADDR 2792
			"00000000000000000000000000000000" , -- ADDR 2793
			"00000000000000000000000000000000" , -- ADDR 2794
			"00000000000000000000000000000000" , -- ADDR 2795
			"00000000000000000000000000000000" , -- ADDR 2796
			"00000000000000000000000000000000" , -- ADDR 2797
			"00000000000000000000000000000000" , -- ADDR 2798
			"00000000000000000000000000000000" , -- ADDR 2799
			"00000000000000000000000000000000" , -- ADDR 2800
			"00000000000000000000000000000000" , -- ADDR 2801
			"00000000000000000000000000000000" , -- ADDR 2802
			"00000000000000000000000000000000" , -- ADDR 2803
			"00000000000000000000000000000000" , -- ADDR 2804
			"00000000000000000000000000000000" , -- ADDR 2805
			"00000000000000000000000000000000" , -- ADDR 2806
			"00000000000000000000000000000000" , -- ADDR 2807
			"00000000000000000000000000000000" , -- ADDR 2808
			"00000000000000000000000000000000" , -- ADDR 2809
			"00000000000000000000000000000000" , -- ADDR 2810
			"00000000000000000000000000000000" , -- ADDR 2811
			"00000000000000000000000000000000" , -- ADDR 2812
			"00000000000000000000000000000000" , -- ADDR 2813
			"00000000000000000000000000000000" , -- ADDR 2814
			"00000000000000000000000000000000" , -- ADDR 2815
			"00000000000000000000000000000000" , -- ADDR 2816
			"00000000000000000000000000000000" , -- ADDR 2817
			"00000000000000000000000000000000" , -- ADDR 2818
			"00000000000000000000000000000000" , -- ADDR 2819
			"00000000000000000000000000000000" , -- ADDR 2820
			"00000000000000000000000000000000" , -- ADDR 2821
			"00000000000000000000000000000000" , -- ADDR 2822
			"00000000000000000000000000000000" , -- ADDR 2823
			"00000000000000000000000000000000" , -- ADDR 2824
			"00000000000000000000000000000000" , -- ADDR 2825
			"00000000000000000000000000000000" , -- ADDR 2826
			"00000000000000000000000000000000" , -- ADDR 2827
			"00000000000000000000000000000000" , -- ADDR 2828
			"00000000000000000000000000000000" , -- ADDR 2829
			"00000000000000000000000000000000" , -- ADDR 2830
			"00000000000000000000000000000000" , -- ADDR 2831
			"00000000000000000000000000000000" , -- ADDR 2832
			"00000000000000000000000000000000" , -- ADDR 2833
			"00000000000000000000000000000000" , -- ADDR 2834
			"00000000000000000000000000000000" , -- ADDR 2835
			"00000000000000000000000000000000" , -- ADDR 2836
			"00000000000000000000000000000000" , -- ADDR 2837
			"00000000000000000000000000000000" , -- ADDR 2838
			"00000000000000000000000000000000" , -- ADDR 2839
			"00000000000000000000000000000000" , -- ADDR 2840
			"00000000000000000000000000000000" , -- ADDR 2841
			"00000000000000000000000000000000" , -- ADDR 2842
			"00000000000000000000000000000000" , -- ADDR 2843
			"00000000000000000000000000000000" , -- ADDR 2844
			"00000000000000000000000000000000" , -- ADDR 2845
			"00000000000000000000000000000000" , -- ADDR 2846
			"00000000000000000000000000000000" , -- ADDR 2847
			"00000000000000000000000000000000" , -- ADDR 2848
			"00000000000000000000000000000000" , -- ADDR 2849
			"00000000000000000000000000000000" , -- ADDR 2850
			"00000000000000000000000000000000" , -- ADDR 2851
			"00000000000000000000000000000000" , -- ADDR 2852
			"00000000000000000000000000000000" , -- ADDR 2853
			"00000000000000000000000000000000" , -- ADDR 2854
			"00000000000000000000000000000000" , -- ADDR 2855
			"00000000000000000000000000000000" , -- ADDR 2856
			"00000000000000000000000000000000" , -- ADDR 2857
			"00000000000000000000000000000000" , -- ADDR 2858
			"00000000000000000000000000000000" , -- ADDR 2859
			"00000000000000000000000000000000" , -- ADDR 2860
			"00000000000000000000000000000000" , -- ADDR 2861
			"00000000000000000000000000000000" , -- ADDR 2862
			"00000000000000000000000000000000" , -- ADDR 2863
			"00000000000000000000000000000000" , -- ADDR 2864
			"00000000000000000000000000000000" , -- ADDR 2865
			"00000000000000000000000000000000" , -- ADDR 2866
			"00000000000000000000000000000000" , -- ADDR 2867
			"00000000000000000000000000000000" , -- ADDR 2868
			"00000000000000000000000000000000" , -- ADDR 2869
			"00000000000000000000000000000000" , -- ADDR 2870
			"00000000000000000000000000000000" , -- ADDR 2871
			"00000000000000000000000000000000" , -- ADDR 2872
			"00000000000000000000000000000000" , -- ADDR 2873
			"00000000000000000000000000000000" , -- ADDR 2874
			"00000000000000000000000000000000" , -- ADDR 2875
			"00000000000000000000000000000000" , -- ADDR 2876
			"00000000000000000000000000000000" , -- ADDR 2877
			"00000000000000000000000000000000" , -- ADDR 2878
			"00000000000000000000000000000000" , -- ADDR 2879
			"00000000000000000000000000000000" , -- ADDR 2880
			"00000000000000000000000000000000" , -- ADDR 2881
			"00000000000000000000000000000000" , -- ADDR 2882
			"00000000000000000000000000000000" , -- ADDR 2883
			"00000000000000000000000000000000" , -- ADDR 2884
			"00000000000000000000000000000000" , -- ADDR 2885
			"00000000000000000000000000000000" , -- ADDR 2886
			"00000000000000000000000000000000" , -- ADDR 2887
			"00000000000000000000000000000000" , -- ADDR 2888
			"00000000000000000000000000000000" , -- ADDR 2889
			"00000000000000000000000000000000" , -- ADDR 2890
			"00000000000000000000000000000000" , -- ADDR 2891
			"00000000000000000000000000000000" , -- ADDR 2892
			"00000000000000000000000000000000" , -- ADDR 2893
			"00000000000000000000000000000000" , -- ADDR 2894
			"00000000000000000000000000000000" , -- ADDR 2895
			"00000000000000000000000000000000" , -- ADDR 2896
			"00000000000000000000000000000000" , -- ADDR 2897
			"00000000000000000000000000000000" , -- ADDR 2898
			"00000000000000000000000000000000" , -- ADDR 2899
			"00000000000000000000000000000000" , -- ADDR 2900
			"00000000000000000000000000000000" , -- ADDR 2901
			"00000000000000000000000000000000" , -- ADDR 2902
			"00000000000000000000000000000000" , -- ADDR 2903
			"00000000000000000000000000000000" , -- ADDR 2904
			"00000000000000000000000000000000" , -- ADDR 2905
			"00000000000000000000000000000000" , -- ADDR 2906
			"00000000000000000000000000000000" , -- ADDR 2907
			"00000000000000000000000000000000" , -- ADDR 2908
			"00000000000000000000000000000000" , -- ADDR 2909
			"00000000000000000000000000000000" , -- ADDR 2910
			"00000000000000000000000000000000" , -- ADDR 2911
			"00000000000000000000000000000000" , -- ADDR 2912
			"00000000000000000000000000000000" , -- ADDR 2913
			"00000000000000000000000000000000" , -- ADDR 2914
			"00000000000000000000000000000000" , -- ADDR 2915
			"00000000000000000000000000000000" , -- ADDR 2916
			"00000000000000000000000000000000" , -- ADDR 2917
			"00000000000000000000000000000000" , -- ADDR 2918
			"00000000000000000000000000000000" , -- ADDR 2919
			"00000000000000000000000000000000" , -- ADDR 2920
			"00000000000000000000000000000000" , -- ADDR 2921
			"00000000000000000000000000000000" , -- ADDR 2922
			"00000000000000000000000000000000" , -- ADDR 2923
			"00000000000000000000000000000000" , -- ADDR 2924
			"00000000000000000000000000000000" , -- ADDR 2925
			"00000000000000000000000000000000" , -- ADDR 2926
			"00000000000000000000000000000000" , -- ADDR 2927
			"00000000000000000000000000000000" , -- ADDR 2928
			"00000000000000000000000000000000" , -- ADDR 2929
			"00000000000000000000000000000000" , -- ADDR 2930
			"00000000000000000000000000000000" , -- ADDR 2931
			"00000000000000000000000000000000" , -- ADDR 2932
			"00000000000000000000000000000000" , -- ADDR 2933
			"00000000000000000000000000000000" , -- ADDR 2934
			"00000000000000000000000000000000" , -- ADDR 2935
			"00000000000000000000000000000000" , -- ADDR 2936
			"00000000000000000000000000000000" , -- ADDR 2937
			"00000000000000000000000000000000" , -- ADDR 2938
			"00000000000000000000000000000000" , -- ADDR 2939
			"00000000000000000000000000000000" , -- ADDR 2940
			"00000000000000000000000000000000" , -- ADDR 2941
			"00000000000000000000000000000000" , -- ADDR 2942
			"00000000000000000000000000000000" , -- ADDR 2943
			"00000000000000000000000000000000" , -- ADDR 2944
			"00000000000000000000000000000000" , -- ADDR 2945
			"00000000000000000000000000000000" , -- ADDR 2946
			"00000000000000000000000000000000" , -- ADDR 2947
			"00000000000000000000000000000000" , -- ADDR 2948
			"00000000000000000000000000000000" , -- ADDR 2949
			"00000000000000000000000000000000" , -- ADDR 2950
			"00000000000000000000000000000000" , -- ADDR 2951
			"00000000000000000000000000000000" , -- ADDR 2952
			"00000000000000000000000000000000" , -- ADDR 2953
			"00000000000000000000000000000000" , -- ADDR 2954
			"00000000000000000000000000000000" , -- ADDR 2955
			"00000000000000000000000000000000" , -- ADDR 2956
			"00000000000000000000000000000000" , -- ADDR 2957
			"00000000000000000000000000000000" , -- ADDR 2958
			"00000000000000000000000000000000" , -- ADDR 2959
			"00000000000000000000000000000000" , -- ADDR 2960
			"00000000000000000000000000000000" , -- ADDR 2961
			"00000000000000000000000000000000" , -- ADDR 2962
			"00000000000000000000000000000000" , -- ADDR 2963
			"00000000000000000000000000000000" , -- ADDR 2964
			"00000000000000000000000000000000" , -- ADDR 2965
			"00000000000000000000000000000000" , -- ADDR 2966
			"00000000000000000000000000000000" , -- ADDR 2967
			"00000000000000000000000000000000" , -- ADDR 2968
			"00000000000000000000000000000000" , -- ADDR 2969
			"00000000000000000000000000000000" , -- ADDR 2970
			"00000000000000000000000000000000" , -- ADDR 2971
			"00000000000000000000000000000000" , -- ADDR 2972
			"00000000000000000000000000000000" , -- ADDR 2973
			"00000000000000000000000000000000" , -- ADDR 2974
			"00000000000000000000000000000000" , -- ADDR 2975
			"00000000000000000000000000000000" , -- ADDR 2976
			"00000000000000000000000000000000" , -- ADDR 2977
			"00000000000000000000000000000000" , -- ADDR 2978
			"00000000000000000000000000000000" , -- ADDR 2979
			"00000000000000000000000000000000" , -- ADDR 2980
			"00000000000000000000000000000000" , -- ADDR 2981
			"00000000000000000000000000000000" , -- ADDR 2982
			"00000000000000000000000000000000" , -- ADDR 2983
			"00000000000000000000000000000000" , -- ADDR 2984
			"00000000000000000000000000000000" , -- ADDR 2985
			"00000000000000000000000000000000" , -- ADDR 2986
			"00000000000000000000000000000000" , -- ADDR 2987
			"00000000000000000000000000000000" , -- ADDR 2988
			"00000000000000000000000000000000" , -- ADDR 2989
			"00000000000000000000000000000000" , -- ADDR 2990
			"00000000000000000000000000000000" , -- ADDR 2991
			"00000000000000000000000000000000" , -- ADDR 2992
			"00000000000000000000000000000000" , -- ADDR 2993
			"00000000000000000000000000000000" , -- ADDR 2994
			"00000000000000000000000000000000" , -- ADDR 2995
			"00000000000000000000000000000000" , -- ADDR 2996
			"00000000000000000000000000000000" , -- ADDR 2997
			"00000000000000000000000000000000" , -- ADDR 2998
			"00000000000000000000000000000000" , -- ADDR 2999
			"00000000000000000000000000000000" , -- ADDR 3000
			"00000000000000000000000000000000" , -- ADDR 3001
			"00000000000000000000000000000000" , -- ADDR 3002
			"00000000000000000000000000000000" , -- ADDR 3003
			"00000000000000000000000000000000" , -- ADDR 3004
			"00000000000000000000000000000000" , -- ADDR 3005
			"00000000000000000000000000000000" , -- ADDR 3006
			"00000000000000000000000000000000" , -- ADDR 3007
			"00000000000000000000000000000000" , -- ADDR 3008
			"00000000000000000000000000000000" , -- ADDR 3009
			"00000000000000000000000000000000" , -- ADDR 3010
			"00000000000000000000000000000000" , -- ADDR 3011
			"00000000000000000000000000000000" , -- ADDR 3012
			"00000000000000000000000000000000" , -- ADDR 3013
			"00000000000000000000000000000000" , -- ADDR 3014
			"00000000000000000000000000000000" , -- ADDR 3015
			"00000000000000000000000000000000" , -- ADDR 3016
			"00000000000000000000000000000000" , -- ADDR 3017
			"00000000000000000000000000000000" , -- ADDR 3018
			"00000000000000000000000000000000" , -- ADDR 3019
			"00000000000000000000000000000000" , -- ADDR 3020
			"00000000000000000000000000000000" , -- ADDR 3021
			"00000000000000000000000000000000" , -- ADDR 3022
			"00000000000000000000000000000000" , -- ADDR 3023
			"00000000000000000000000000000000" , -- ADDR 3024
			"00000000000000000000000000000000" , -- ADDR 3025
			"00000000000000000000000000000000" , -- ADDR 3026
			"00000000000000000000000000000000" , -- ADDR 3027
			"00000000000000000000000000000000" , -- ADDR 3028
			"00000000000000000000000000000000" , -- ADDR 3029
			"00000000000000000000000000000000" , -- ADDR 3030
			"00000000000000000000000000000000" , -- ADDR 3031
			"00000000000000000000000000000000" , -- ADDR 3032
			"00000000000000000000000000000000" , -- ADDR 3033
			"00000000000000000000000000000000" , -- ADDR 3034
			"00000000000000000000000000000000" , -- ADDR 3035
			"00000000000000000000000000000000" , -- ADDR 3036
			"00000000000000000000000000000000" , -- ADDR 3037
			"00000000000000000000000000000000" , -- ADDR 3038
			"00000000000000000000000000000000" , -- ADDR 3039
			"00000000000000000000000000000000" , -- ADDR 3040
			"00000000000000000000000000000000" , -- ADDR 3041
			"00000000000000000000000000000000" , -- ADDR 3042
			"00000000000000000000000000000000" , -- ADDR 3043
			"00000000000000000000000000000000" , -- ADDR 3044
			"00000000000000000000000000000000" , -- ADDR 3045
			"00000000000000000000000000000000" , -- ADDR 3046
			"00000000000000000000000000000000" , -- ADDR 3047
			"00000000000000000000000000000000" , -- ADDR 3048
			"00000000000000000000000000000000" , -- ADDR 3049
			"00000000000000000000000000000000" , -- ADDR 3050
			"00000000000000000000000000000000" , -- ADDR 3051
			"00000000000000000000000000000000" , -- ADDR 3052
			"00000000000000000000000000000000" , -- ADDR 3053
			"00000000000000000000000000000000" , -- ADDR 3054
			"00000000000000000000000000000000" , -- ADDR 3055
			"00000000000000000000000000000000" , -- ADDR 3056
			"00000000000000000000000000000000" , -- ADDR 3057
			"00000000000000000000000000000000" , -- ADDR 3058
			"00000000000000000000000000000000" , -- ADDR 3059
			"00000000000000000000000000000000" , -- ADDR 3060
			"00000000000000000000000000000000" , -- ADDR 3061
			"00000000000000000000000000000000" , -- ADDR 3062
			"00000000000000000000000000000000" , -- ADDR 3063
			"00000000000000000000000000000000" , -- ADDR 3064
			"00000000000000000000000000000000" , -- ADDR 3065
			"00000000000000000000000000000000" , -- ADDR 3066
			"00000000000000000000000000000000" , -- ADDR 3067
			"00000000000000000000000000000000" , -- ADDR 3068
			"00000000000000000000000000000000" , -- ADDR 3069
			"00000000000000000000000000000000" , -- ADDR 3070
			"00000000000000000000000000000000" , -- ADDR 3071
			"00000000000000000000000000000000" , -- ADDR 3072
			"00000000000000000000000000000000" , -- ADDR 3073
			"00000000000000000000000000000000" , -- ADDR 3074
			"00000000000000000000000000000000" , -- ADDR 3075
			"00000000000000000000000000000000" , -- ADDR 3076
			"00000000000000000000000000000000" , -- ADDR 3077
			"00000000000000000000000000000000" , -- ADDR 3078
			"00000000000000000000000000000000" , -- ADDR 3079
			"00000000000000000000000000000000" , -- ADDR 3080
			"00000000000000000000000000000000" , -- ADDR 3081
			"00000000000000000000000000000000" , -- ADDR 3082
			"00000000000000000000000000000000" , -- ADDR 3083
			"00000000000000000000000000000000" , -- ADDR 3084
			"00000000000000000000000000000000" , -- ADDR 3085
			"00000000000000000000000000000000" , -- ADDR 3086
			"00000000000000000000000000000000" , -- ADDR 3087
			"00000000000000000000000000000000" , -- ADDR 3088
			"00000000000000000000000000000000" , -- ADDR 3089
			"00000000000000000000000000000000" , -- ADDR 3090
			"00000000000000000000000000000000" , -- ADDR 3091
			"00000000000000000000000000000000" , -- ADDR 3092
			"00000000000000000000000000000000" , -- ADDR 3093
			"00000000000000000000000000000000" , -- ADDR 3094
			"00000000000000000000000000000000" , -- ADDR 3095
			"00000000000000000000000000000000" , -- ADDR 3096
			"00000000000000000000000000000000" , -- ADDR 3097
			"00000000000000000000000000000000" , -- ADDR 3098
			"00000000000000000000000000000000" , -- ADDR 3099
			"00000000000000000000000000000000" , -- ADDR 3100
			"00000000000000000000000000000000" , -- ADDR 3101
			"00000000000000000000000000000000" , -- ADDR 3102
			"00000000000000000000000000000000" , -- ADDR 3103
			"00000000000000000000000000000000" , -- ADDR 3104
			"00000000000000000000000000000000" , -- ADDR 3105
			"00000000000000000000000000000000" , -- ADDR 3106
			"00000000000000000000000000000000" , -- ADDR 3107
			"00000000000000000000000000000000" , -- ADDR 3108
			"00000000000000000000000000000000" , -- ADDR 3109
			"00000000000000000000000000000000" , -- ADDR 3110
			"00000000000000000000000000000000" , -- ADDR 3111
			"00000000000000000000000000000000" , -- ADDR 3112
			"00000000000000000000000000000000" , -- ADDR 3113
			"00000000000000000000000000000000" , -- ADDR 3114
			"00000000000000000000000000000000" , -- ADDR 3115
			"00000000000000000000000000000000" , -- ADDR 3116
			"00000000000000000000000000000000" , -- ADDR 3117
			"00000000000000000000000000000000" , -- ADDR 3118
			"00000000000000000000000000000000" , -- ADDR 3119
			"00000000000000000000000000000000" , -- ADDR 3120
			"00000000000000000000000000000000" , -- ADDR 3121
			"00000000000000000000000000000000" , -- ADDR 3122
			"00000000000000000000000000000000" , -- ADDR 3123
			"00000000000000000000000000000000" , -- ADDR 3124
			"00000000000000000000000000000000" , -- ADDR 3125
			"00000000000000000000000000000000" , -- ADDR 3126
			"00000000000000000000000000000000" , -- ADDR 3127
			"00000000000000000000000000000000" , -- ADDR 3128
			"00000000000000000000000000000000" , -- ADDR 3129
			"00000000000000000000000000000000" , -- ADDR 3130
			"00000000000000000000000000000000" , -- ADDR 3131
			"00000000000000000000000000000000" , -- ADDR 3132
			"00000000000000000000000000000000" , -- ADDR 3133
			"00000000000000000000000000000000" , -- ADDR 3134
			"00000000000000000000000000000000" , -- ADDR 3135
			"00000000000000000000000000000000" , -- ADDR 3136
			"00000000000000000000000000000000" , -- ADDR 3137
			"00000000000000000000000000000000" , -- ADDR 3138
			"00000000000000000000000000000000" , -- ADDR 3139
			"00000000000000000000000000000000" , -- ADDR 3140
			"00000000000000000000000000000000" , -- ADDR 3141
			"00000000000000000000000000000000" , -- ADDR 3142
			"00000000000000000000000000000000" , -- ADDR 3143
			"00000000000000000000000000000000" , -- ADDR 3144
			"00000000000000000000000000000000" , -- ADDR 3145
			"00000000000000000000000000000000" , -- ADDR 3146
			"00000000000000000000000000000000" , -- ADDR 3147
			"00000000000000000000000000000000" , -- ADDR 3148
			"00000000000000000000000000000000" , -- ADDR 3149
			"00000000000000000000000000000000" , -- ADDR 3150
			"00000000000000000000000000000000" , -- ADDR 3151
			"00000000000000000000000000000000" , -- ADDR 3152
			"00000000000000000000000000000000" , -- ADDR 3153
			"00000000000000000000000000000000" , -- ADDR 3154
			"00000000000000000000000000000000" , -- ADDR 3155
			"00000000000000000000000000000000" , -- ADDR 3156
			"00000000000000000000000000000000" , -- ADDR 3157
			"00000000000000000000000000000000" , -- ADDR 3158
			"00000000000000000000000000000000" , -- ADDR 3159
			"00000000000000000000000000000000" , -- ADDR 3160
			"00000000000000000000000000000000" , -- ADDR 3161
			"00000000000000000000000000000000" , -- ADDR 3162
			"00000000000000000000000000000000" , -- ADDR 3163
			"00000000000000000000000000000000" , -- ADDR 3164
			"00000000000000000000000000000000" , -- ADDR 3165
			"00000000000000000000000000000000" , -- ADDR 3166
			"00000000000000000000000000000000" , -- ADDR 3167
			"00000000000000000000000000000000" , -- ADDR 3168
			"00000000000000000000000000000000" , -- ADDR 3169
			"00000000000000000000000000000000" , -- ADDR 3170
			"00000000000000000000000000000000" , -- ADDR 3171
			"00000000000000000000000000000000" , -- ADDR 3172
			"00000000000000000000000000000000" , -- ADDR 3173
			"00000000000000000000000000000000" , -- ADDR 3174
			"00000000000000000000000000000000" , -- ADDR 3175
			"00000000000000000000000000000000" , -- ADDR 3176
			"00000000000000000000000000000000" , -- ADDR 3177
			"00000000000000000000000000000000" , -- ADDR 3178
			"00000000000000000000000000000000" , -- ADDR 3179
			"00000000000000000000000000000000" , -- ADDR 3180
			"00000000000000000000000000000000" , -- ADDR 3181
			"00000000000000000000000000000000" , -- ADDR 3182
			"00000000000000000000000000000000" , -- ADDR 3183
			"00000000000000000000000000000000" , -- ADDR 3184
			"00000000000000000000000000000000" , -- ADDR 3185
			"00000000000000000000000000000000" , -- ADDR 3186
			"00000000000000000000000000000000" , -- ADDR 3187
			"00000000000000000000000000000000" , -- ADDR 3188
			"00000000000000000000000000000000" , -- ADDR 3189
			"00000000000000000000000000000000" , -- ADDR 3190
			"00000000000000000000000000000000" , -- ADDR 3191
			"00000000000000000000000000000000" , -- ADDR 3192
			"00000000000000000000000000000000" , -- ADDR 3193
			"00000000000000000000000000000000" , -- ADDR 3194
			"00000000000000000000000000000000" , -- ADDR 3195
			"00000000000000000000000000000000" , -- ADDR 3196
			"00000000000000000000000000000000" , -- ADDR 3197
			"00000000000000000000000000000000" , -- ADDR 3198
			"00000000000000000000000000000000" , -- ADDR 3199
			"00000000000000000000000000000000" , -- ADDR 3200
			"00000000000000000000000000000000" , -- ADDR 3201
			"00000000000000000000000000000000" , -- ADDR 3202
			"00000000000000000000000000000000" , -- ADDR 3203
			"00000000000000000000000000000000" , -- ADDR 3204
			"00000000000000000000000000000000" , -- ADDR 3205
			"00000000000000000000000000000000" , -- ADDR 3206
			"00000000000000000000000000000000" , -- ADDR 3207
			"00000000000000000000000000000000" , -- ADDR 3208
			"00000000000000000000000000000000" , -- ADDR 3209
			"00000000000000000000000000000000" , -- ADDR 3210
			"00000000000000000000000000000000" , -- ADDR 3211
			"00000000000000000000000000000000" , -- ADDR 3212
			"00000000000000000000000000000000" , -- ADDR 3213
			"00000000000000000000000000000000" , -- ADDR 3214
			"00000000000000000000000000000000" , -- ADDR 3215
			"00000000000000000000000000000000" , -- ADDR 3216
			"00000000000000000000000000000000" , -- ADDR 3217
			"00000000000000000000000000000000" , -- ADDR 3218
			"00000000000000000000000000000000" , -- ADDR 3219
			"00000000000000000000000000000000" , -- ADDR 3220
			"00000000000000000000000000000000" , -- ADDR 3221
			"00000000000000000000000000000000" , -- ADDR 3222
			"00000000000000000000000000000000" , -- ADDR 3223
			"00000000000000000000000000000000" , -- ADDR 3224
			"00000000000000000000000000000000" , -- ADDR 3225
			"00000000000000000000000000000000" , -- ADDR 3226
			"00000000000000000000000000000000" , -- ADDR 3227
			"00000000000000000000000000000000" , -- ADDR 3228
			"00000000000000000000000000000000" , -- ADDR 3229
			"00000000000000000000000000000000" , -- ADDR 3230
			"00000000000000000000000000000000" , -- ADDR 3231
			"00000000000000000000000000000000" , -- ADDR 3232
			"00000000000000000000000000000000" , -- ADDR 3233
			"00000000000000000000000000000000" , -- ADDR 3234
			"00000000000000000000000000000000" , -- ADDR 3235
			"00000000000000000000000000000000" , -- ADDR 3236
			"00000000000000000000000000000000" , -- ADDR 3237
			"00000000000000000000000000000000" , -- ADDR 3238
			"00000000000000000000000000000000" , -- ADDR 3239
			"00000000000000000000000000000000" , -- ADDR 3240
			"00000000000000000000000000000000" , -- ADDR 3241
			"00000000000000000000000000000000" , -- ADDR 3242
			"00000000000000000000000000000000" , -- ADDR 3243
			"00000000000000000000000000000000" , -- ADDR 3244
			"00000000000000000000000000000000" , -- ADDR 3245
			"00000000000000000000000000000000" , -- ADDR 3246
			"00000000000000000000000000000000" , -- ADDR 3247
			"00000000000000000000000000000000" , -- ADDR 3248
			"00000000000000000000000000000000" , -- ADDR 3249
			"00000000000000000000000000000000" , -- ADDR 3250
			"00000000000000000000000000000000" , -- ADDR 3251
			"00000000000000000000000000000000" , -- ADDR 3252
			"00000000000000000000000000000000" , -- ADDR 3253
			"00000000000000000000000000000000" , -- ADDR 3254
			"00000000000000000000000000000000" , -- ADDR 3255
			"00000000000000000000000000000000" , -- ADDR 3256
			"00000000000000000000000000000000" , -- ADDR 3257
			"00000000000000000000000000000000" , -- ADDR 3258
			"00000000000000000000000000000000" , -- ADDR 3259
			"00000000000000000000000000000000" , -- ADDR 3260
			"00000000000000000000000000000000" , -- ADDR 3261
			"00000000000000000000000000000000" , -- ADDR 3262
			"00000000000000000000000000000000" , -- ADDR 3263
			"00000000000000000000000000000000" , -- ADDR 3264
			"00000000000000000000000000000000" , -- ADDR 3265
			"00000000000000000000000000000000" , -- ADDR 3266
			"00000000000000000000000000000000" , -- ADDR 3267
			"00000000000000000000000000000000" , -- ADDR 3268
			"00000000000000000000000000000000" , -- ADDR 3269
			"00000000000000000000000000000000" , -- ADDR 3270
			"00000000000000000000000000000000" , -- ADDR 3271
			"00000000000000000000000000000000" , -- ADDR 3272
			"00000000000000000000000000000000" , -- ADDR 3273
			"00000000000000000000000000000000" , -- ADDR 3274
			"00000000000000000000000000000000" , -- ADDR 3275
			"00000000000000000000000000000000" , -- ADDR 3276
			"00000000000000000000000000000000" , -- ADDR 3277
			"00000000000000000000000000000000" , -- ADDR 3278
			"00000000000000000000000000000000" , -- ADDR 3279
			"00000000000000000000000000000000" , -- ADDR 3280
			"00000000000000000000000000000000" , -- ADDR 3281
			"00000000000000000000000000000000" , -- ADDR 3282
			"00000000000000000000000000000000" , -- ADDR 3283
			"00000000000000000000000000000000" , -- ADDR 3284
			"00000000000000000000000000000000" , -- ADDR 3285
			"00000000000000000000000000000000" , -- ADDR 3286
			"00000000000000000000000000000000" , -- ADDR 3287
			"00000000000000000000000000000000" , -- ADDR 3288
			"00000000000000000000000000000000" , -- ADDR 3289
			"00000000000000000000000000000000" , -- ADDR 3290
			"00000000000000000000000000000000" , -- ADDR 3291
			"00000000000000000000000000000000" , -- ADDR 3292
			"00000000000000000000000000000000" , -- ADDR 3293
			"00000000000000000000000000000000" , -- ADDR 3294
			"00000000000000000000000000000000" , -- ADDR 3295
			"00000000000000000000000000000000" , -- ADDR 3296
			"00000000000000000000000000000000" , -- ADDR 3297
			"00000000000000000000000000000000" , -- ADDR 3298
			"00000000000000000000000000000000" , -- ADDR 3299
			"00000000000000000000000000000000" , -- ADDR 3300
			"00000000000000000000000000000000" , -- ADDR 3301
			"00000000000000000000000000000000" , -- ADDR 3302
			"00000000000000000000000000000000" , -- ADDR 3303
			"00000000000000000000000000000000" , -- ADDR 3304
			"00000000000000000000000000000000" , -- ADDR 3305
			"00000000000000000000000000000000" , -- ADDR 3306
			"00000000000000000000000000000000" , -- ADDR 3307
			"00000000000000000000000000000000" , -- ADDR 3308
			"00000000000000000000000000000000" , -- ADDR 3309
			"00000000000000000000000000000000" , -- ADDR 3310
			"00000000000000000000000000000000" , -- ADDR 3311
			"00000000000000000000000000000000" , -- ADDR 3312
			"00000000000000000000000000000000" , -- ADDR 3313
			"00000000000000000000000000000000" , -- ADDR 3314
			"00000000000000000000000000000000" , -- ADDR 3315
			"00000000000000000000000000000000" , -- ADDR 3316
			"00000000000000000000000000000000" , -- ADDR 3317
			"00000000000000000000000000000000" , -- ADDR 3318
			"00000000000000000000000000000000" , -- ADDR 3319
			"00000000000000000000000000000000" , -- ADDR 3320
			"00000000000000000000000000000000" , -- ADDR 3321
			"00000000000000000000000000000000" , -- ADDR 3322
			"00000000000000000000000000000000" , -- ADDR 3323
			"00000000000000000000000000000000" , -- ADDR 3324
			"00000000000000000000000000000000" , -- ADDR 3325
			"00000000000000000000000000000000" , -- ADDR 3326
			"00000000000000000000000000000000" , -- ADDR 3327
			"00000000000000000000000000000000" , -- ADDR 3328
			"00000000000000000000000000000000" , -- ADDR 3329
			"00000000000000000000000000000000" , -- ADDR 3330
			"00000000000000000000000000000000" , -- ADDR 3331
			"00000000000000000000000000000000" , -- ADDR 3332
			"00000000000000000000000000000000" , -- ADDR 3333
			"00000000000000000000000000000000" , -- ADDR 3334
			"00000000000000000000000000000000" , -- ADDR 3335
			"00000000000000000000000000000000" , -- ADDR 3336
			"00000000000000000000000000000000" , -- ADDR 3337
			"00000000000000000000000000000000" , -- ADDR 3338
			"00000000000000000000000000000000" , -- ADDR 3339
			"00000000000000000000000000000000" , -- ADDR 3340
			"00000000000000000000000000000000" , -- ADDR 3341
			"00000000000000000000000000000000" , -- ADDR 3342
			"00000000000000000000000000000000" , -- ADDR 3343
			"00000000000000000000000000000000" , -- ADDR 3344
			"00000000000000000000000000000000" , -- ADDR 3345
			"00000000000000000000000000000000" , -- ADDR 3346
			"00000000000000000000000000000000" , -- ADDR 3347
			"00000000000000000000000000000000" , -- ADDR 3348
			"00000000000000000000000000000000" , -- ADDR 3349
			"00000000000000000000000000000000" , -- ADDR 3350
			"00000000000000000000000000000000" , -- ADDR 3351
			"00000000000000000000000000000000" , -- ADDR 3352
			"00000000000000000000000000000000" , -- ADDR 3353
			"00000000000000000000000000000000" , -- ADDR 3354
			"00000000000000000000000000000000" , -- ADDR 3355
			"00000000000000000000000000000000" , -- ADDR 3356
			"00000000000000000000000000000000" , -- ADDR 3357
			"00000000000000000000000000000000" , -- ADDR 3358
			"00000000000000000000000000000000" , -- ADDR 3359
			"00000000000000000000000000000000" , -- ADDR 3360
			"00000000000000000000000000000000" , -- ADDR 3361
			"00000000000000000000000000000000" , -- ADDR 3362
			"00000000000000000000000000000000" , -- ADDR 3363
			"00000000000000000000000000000000" , -- ADDR 3364
			"00000000000000000000000000000000" , -- ADDR 3365
			"00000000000000000000000000000000" , -- ADDR 3366
			"00000000000000000000000000000000" , -- ADDR 3367
			"00000000000000000000000000000000" , -- ADDR 3368
			"00000000000000000000000000000000" , -- ADDR 3369
			"00000000000000000000000000000000" , -- ADDR 3370
			"00000000000000000000000000000000" , -- ADDR 3371
			"00000000000000000000000000000000" , -- ADDR 3372
			"00000000000000000000000000000000" , -- ADDR 3373
			"00000000000000000000000000000000" , -- ADDR 3374
			"00000000000000000000000000000000" , -- ADDR 3375
			"00000000000000000000000000000000" , -- ADDR 3376
			"00000000000000000000000000000000" , -- ADDR 3377
			"00000000000000000000000000000000" , -- ADDR 3378
			"00000000000000000000000000000000" , -- ADDR 3379
			"00000000000000000000000000000000" , -- ADDR 3380
			"00000000000000000000000000000000" , -- ADDR 3381
			"00000000000000000000000000000000" , -- ADDR 3382
			"00000000000000000000000000000000" , -- ADDR 3383
			"00000000000000000000000000000000" , -- ADDR 3384
			"00000000000000000000000000000000" , -- ADDR 3385
			"00000000000000000000000000000000" , -- ADDR 3386
			"00000000000000000000000000000000" , -- ADDR 3387
			"00000000000000000000000000000000" , -- ADDR 3388
			"00000000000000000000000000000000" , -- ADDR 3389
			"00000000000000000000000000000000" , -- ADDR 3390
			"00000000000000000000000000000000" , -- ADDR 3391
			"00000000000000000000000000000000" , -- ADDR 3392
			"00000000000000000000000000000000" , -- ADDR 3393
			"00000000000000000000000000000000" , -- ADDR 3394
			"00000000000000000000000000000000" , -- ADDR 3395
			"00000000000000000000000000000000" , -- ADDR 3396
			"00000000000000000000000000000000" , -- ADDR 3397
			"00000000000000000000000000000000" , -- ADDR 3398
			"00000000000000000000000000000000" , -- ADDR 3399
			"00000000000000000000000000000000" , -- ADDR 3400
			"00000000000000000000000000000000" , -- ADDR 3401
			"00000000000000000000000000000000" , -- ADDR 3402
			"00000000000000000000000000000000" , -- ADDR 3403
			"00000000000000000000000000000000" , -- ADDR 3404
			"00000000000000000000000000000000" , -- ADDR 3405
			"00000000000000000000000000000000" , -- ADDR 3406
			"00000000000000000000000000000000" , -- ADDR 3407
			"00000000000000000000000000000000" , -- ADDR 3408
			"00000000000000000000000000000000" , -- ADDR 3409
			"00000000000000000000000000000000" , -- ADDR 3410
			"00000000000000000000000000000000" , -- ADDR 3411
			"00000000000000000000000000000000" , -- ADDR 3412
			"00000000000000000000000000000000" , -- ADDR 3413
			"00000000000000000000000000000000" , -- ADDR 3414
			"00000000000000000000000000000000" , -- ADDR 3415
			"00000000000000000000000000000000" , -- ADDR 3416
			"00000000000000000000000000000000" , -- ADDR 3417
			"00000000000000000000000000000000" , -- ADDR 3418
			"00000000000000000000000000000000" , -- ADDR 3419
			"00000000000000000000000000000000" , -- ADDR 3420
			"00000000000000000000000000000000" , -- ADDR 3421
			"00000000000000000000000000000000" , -- ADDR 3422
			"00000000000000000000000000000000" , -- ADDR 3423
			"00000000000000000000000000000000" , -- ADDR 3424
			"00000000000000000000000000000000" , -- ADDR 3425
			"00000000000000000000000000000000" , -- ADDR 3426
			"00000000000000000000000000000000" , -- ADDR 3427
			"00000000000000000000000000000000" , -- ADDR 3428
			"00000000000000000000000000000000" , -- ADDR 3429
			"00000000000000000000000000000000" , -- ADDR 3430
			"00000000000000000000000000000000" , -- ADDR 3431
			"00000000000000000000000000000000" , -- ADDR 3432
			"00000000000000000000000000000000" , -- ADDR 3433
			"00000000000000000000000000000000" , -- ADDR 3434
			"00000000000000000000000000000000" , -- ADDR 3435
			"00000000000000000000000000000000" , -- ADDR 3436
			"00000000000000000000000000000000" , -- ADDR 3437
			"00000000000000000000000000000000" , -- ADDR 3438
			"00000000000000000000000000000000" , -- ADDR 3439
			"00000000000000000000000000000000" , -- ADDR 3440
			"00000000000000000000000000000000" , -- ADDR 3441
			"00000000000000000000000000000000" , -- ADDR 3442
			"00000000000000000000000000000000" , -- ADDR 3443
			"00000000000000000000000000000000" , -- ADDR 3444
			"00000000000000000000000000000000" , -- ADDR 3445
			"00000000000000000000000000000000" , -- ADDR 3446
			"00000000000000000000000000000000" , -- ADDR 3447
			"00000000000000000000000000000000" , -- ADDR 3448
			"00000000000000000000000000000000" , -- ADDR 3449
			"00000000000000000000000000000000" , -- ADDR 3450
			"00000000000000000000000000000000" , -- ADDR 3451
			"00000000000000000000000000000000" , -- ADDR 3452
			"00000000000000000000000000000000" , -- ADDR 3453
			"00000000000000000000000000000000" , -- ADDR 3454
			"00000000000000000000000000000000" , -- ADDR 3455
			"00000000000000000000000000000000" , -- ADDR 3456
			"00000000000000000000000000000000" , -- ADDR 3457
			"00000000000000000000000000000000" , -- ADDR 3458
			"00000000000000000000000000000000" , -- ADDR 3459
			"00000000000000000000000000000000" , -- ADDR 3460
			"00000000000000000000000000000000" , -- ADDR 3461
			"00000000000000000000000000000000" , -- ADDR 3462
			"00000000000000000000000000000000" , -- ADDR 3463
			"00000000000000000000000000000000" , -- ADDR 3464
			"00000000000000000000000000000000" , -- ADDR 3465
			"00000000000000000000000000000000" , -- ADDR 3466
			"00000000000000000000000000000000" , -- ADDR 3467
			"00000000000000000000000000000000" , -- ADDR 3468
			"00000000000000000000000000000000" , -- ADDR 3469
			"00000000000000000000000000000000" , -- ADDR 3470
			"00000000000000000000000000000000" , -- ADDR 3471
			"00000000000000000000000000000000" , -- ADDR 3472
			"00000000000000000000000000000000" , -- ADDR 3473
			"00000000000000000000000000000000" , -- ADDR 3474
			"00000000000000000000000000000000" , -- ADDR 3475
			"00000000000000000000000000000000" , -- ADDR 3476
			"00000000000000000000000000000000" , -- ADDR 3477
			"00000000000000000000000000000000" , -- ADDR 3478
			"00000000000000000000000000000000" , -- ADDR 3479
			"00000000000000000000000000000000" , -- ADDR 3480
			"00000000000000000000000000000000" , -- ADDR 3481
			"00000000000000000000000000000000" , -- ADDR 3482
			"00000000000000000000000000000000" , -- ADDR 3483
			"00000000000000000000000000000000" , -- ADDR 3484
			"00000000000000000000000000000000" , -- ADDR 3485
			"00000000000000000000000000000000" , -- ADDR 3486
			"00000000000000000000000000000000" , -- ADDR 3487
			"00000000000000000000000000000000" , -- ADDR 3488
			"00000000000000000000000000000000" , -- ADDR 3489
			"00000000000000000000000000000000" , -- ADDR 3490
			"00000000000000000000000000000000" , -- ADDR 3491
			"00000000000000000000000000000000" , -- ADDR 3492
			"00000000000000000000000000000000" , -- ADDR 3493
			"00000000000000000000000000000000" , -- ADDR 3494
			"00000000000000000000000000000000" , -- ADDR 3495
			"00000000000000000000000000000000" , -- ADDR 3496
			"00000000000000000000000000000000" , -- ADDR 3497
			"00000000000000000000000000000000" , -- ADDR 3498
			"00000000000000000000000000000000" , -- ADDR 3499
			"00000000000000000000000000000000" , -- ADDR 3500
			"00000000000000000000000000000000" , -- ADDR 3501
			"00000000000000000000000000000000" , -- ADDR 3502
			"00000000000000000000000000000000" , -- ADDR 3503
			"00000000000000000000000000000000" , -- ADDR 3504
			"00000000000000000000000000000000" , -- ADDR 3505
			"00000000000000000000000000000000" , -- ADDR 3506
			"00000000000000000000000000000000" , -- ADDR 3507
			"00000000000000000000000000000000" , -- ADDR 3508
			"00000000000000000000000000000000" , -- ADDR 3509
			"00000000000000000000000000000000" , -- ADDR 3510
			"00000000000000000000000000000000" , -- ADDR 3511
			"00000000000000000000000000000000" , -- ADDR 3512
			"00000000000000000000000000000000" , -- ADDR 3513
			"00000000000000000000000000000000" , -- ADDR 3514
			"00000000000000000000000000000000" , -- ADDR 3515
			"00000000000000000000000000000000" , -- ADDR 3516
			"00000000000000000000000000000000" , -- ADDR 3517
			"00000000000000000000000000000000" , -- ADDR 3518
			"00000000000000000000000000000000" , -- ADDR 3519
			"00000000000000000000000000000000" , -- ADDR 3520
			"00000000000000000000000000000000" , -- ADDR 3521
			"00000000000000000000000000000000" , -- ADDR 3522
			"00000000000000000000000000000000" , -- ADDR 3523
			"00000000000000000000000000000000" , -- ADDR 3524
			"00000000000000000000000000000000" , -- ADDR 3525
			"00000000000000000000000000000000" , -- ADDR 3526
			"00000000000000000000000000000000" , -- ADDR 3527
			"00000000000000000000000000000000" , -- ADDR 3528
			"00000000000000000000000000000000" , -- ADDR 3529
			"00000000000000000000000000000000" , -- ADDR 3530
			"00000000000000000000000000000000" , -- ADDR 3531
			"00000000000000000000000000000000" , -- ADDR 3532
			"00000000000000000000000000000000" , -- ADDR 3533
			"00000000000000000000000000000000" , -- ADDR 3534
			"00000000000000000000000000000000" , -- ADDR 3535
			"00000000000000000000000000000000" , -- ADDR 3536
			"00000000000000000000000000000000" , -- ADDR 3537
			"00000000000000000000000000000000" , -- ADDR 3538
			"00000000000000000000000000000000" , -- ADDR 3539
			"00000000000000000000000000000000" , -- ADDR 3540
			"00000000000000000000000000000000" , -- ADDR 3541
			"00000000000000000000000000000000" , -- ADDR 3542
			"00000000000000000000000000000000" , -- ADDR 3543
			"00000000000000000000000000000000" , -- ADDR 3544
			"00000000000000000000000000000000" , -- ADDR 3545
			"00000000000000000000000000000000" , -- ADDR 3546
			"00000000000000000000000000000000" , -- ADDR 3547
			"00000000000000000000000000000000" , -- ADDR 3548
			"00000000000000000000000000000000" , -- ADDR 3549
			"00000000000000000000000000000000" , -- ADDR 3550
			"00000000000000000000000000000000" , -- ADDR 3551
			"00000000000000000000000000000000" , -- ADDR 3552
			"00000000000000000000000000000000" , -- ADDR 3553
			"00000000000000000000000000000000" , -- ADDR 3554
			"00000000000000000000000000000000" , -- ADDR 3555
			"00000000000000000000000000000000" , -- ADDR 3556
			"00000000000000000000000000000000" , -- ADDR 3557
			"00000000000000000000000000000000" , -- ADDR 3558
			"00000000000000000000000000000000" , -- ADDR 3559
			"00000000000000000000000000000000" , -- ADDR 3560
			"00000000000000000000000000000000" , -- ADDR 3561
			"00000000000000000000000000000000" , -- ADDR 3562
			"00000000000000000000000000000000" , -- ADDR 3563
			"00000000000000000000000000000000" , -- ADDR 3564
			"00000000000000000000000000000000" , -- ADDR 3565
			"00000000000000000000000000000000" , -- ADDR 3566
			"00000000000000000000000000000000" , -- ADDR 3567
			"00000000000000000000000000000000" , -- ADDR 3568
			"00000000000000000000000000000000" , -- ADDR 3569
			"00000000000000000000000000000000" , -- ADDR 3570
			"00000000000000000000000000000000" , -- ADDR 3571
			"00000000000000000000000000000000" , -- ADDR 3572
			"00000000000000000000000000000000" , -- ADDR 3573
			"00000000000000000000000000000000" , -- ADDR 3574
			"00000000000000000000000000000000" , -- ADDR 3575
			"00000000000000000000000000000000" , -- ADDR 3576
			"00000000000000000000000000000000" , -- ADDR 3577
			"00000000000000000000000000000000" , -- ADDR 3578
			"00000000000000000000000000000000" , -- ADDR 3579
			"00000000000000000000000000000000" , -- ADDR 3580
			"00000000000000000000000000000000" , -- ADDR 3581
			"00000000000000000000000000000000" , -- ADDR 3582
			"00000000000000000000000000000000" , -- ADDR 3583
			"00000000000000000000000000000000" , -- ADDR 3584
			"00000000000000000000000000000000" , -- ADDR 3585
			"00000000000000000000000000000000" , -- ADDR 3586
			"00000000000000000000000000000000" , -- ADDR 3587
			"00000000000000000000000000000000" , -- ADDR 3588
			"00000000000000000000000000000000" , -- ADDR 3589
			"00000000000000000000000000000000" , -- ADDR 3590
			"00000000000000000000000000000000" , -- ADDR 3591
			"00000000000000000000000000000000" , -- ADDR 3592
			"00000000000000000000000000000000" , -- ADDR 3593
			"00000000000000000000000000000000" , -- ADDR 3594
			"00000000000000000000000000000000" , -- ADDR 3595
			"00000000000000000000000000000000" , -- ADDR 3596
			"00000000000000000000000000000000" , -- ADDR 3597
			"00000000000000000000000000000000" , -- ADDR 3598
			"00000000000000000000000000000000" , -- ADDR 3599
			"00000000000000000000000000000000" , -- ADDR 3600
			"00000000000000000000000000000000" , -- ADDR 3601
			"00000000000000000000000000000000" , -- ADDR 3602
			"00000000000000000000000000000000" , -- ADDR 3603
			"00000000000000000000000000000000" , -- ADDR 3604
			"00000000000000000000000000000000" , -- ADDR 3605
			"00000000000000000000000000000000" , -- ADDR 3606
			"00000000000000000000000000000000" , -- ADDR 3607
			"00000000000000000000000000000000" , -- ADDR 3608
			"00000000000000000000000000000000" , -- ADDR 3609
			"00000000000000000000000000000000" , -- ADDR 3610
			"00000000000000000000000000000000" , -- ADDR 3611
			"00000000000000000000000000000000" , -- ADDR 3612
			"00000000000000000000000000000000" , -- ADDR 3613
			"00000000000000000000000000000000" , -- ADDR 3614
			"00000000000000000000000000000000" , -- ADDR 3615
			"00000000000000000000000000000000" , -- ADDR 3616
			"00000000000000000000000000000000" , -- ADDR 3617
			"00000000000000000000000000000000" , -- ADDR 3618
			"00000000000000000000000000000000" , -- ADDR 3619
			"00000000000000000000000000000000" , -- ADDR 3620
			"00000000000000000000000000000000" , -- ADDR 3621
			"00000000000000000000000000000000" , -- ADDR 3622
			"00000000000000000000000000000000" , -- ADDR 3623
			"00000000000000000000000000000000" , -- ADDR 3624
			"00000000000000000000000000000000" , -- ADDR 3625
			"00000000000000000000000000000000" , -- ADDR 3626
			"00000000000000000000000000000000" , -- ADDR 3627
			"00000000000000000000000000000000" , -- ADDR 3628
			"00000000000000000000000000000000" , -- ADDR 3629
			"00000000000000000000000000000000" , -- ADDR 3630
			"00000000000000000000000000000000" , -- ADDR 3631
			"00000000000000000000000000000000" , -- ADDR 3632
			"00000000000000000000000000000000" , -- ADDR 3633
			"00000000000000000000000000000000" , -- ADDR 3634
			"00000000000000000000000000000000" , -- ADDR 3635
			"00000000000000000000000000000000" , -- ADDR 3636
			"00000000000000000000000000000000" , -- ADDR 3637
			"00000000000000000000000000000000" , -- ADDR 3638
			"00000000000000000000000000000000" , -- ADDR 3639
			"00000000000000000000000000000000" , -- ADDR 3640
			"00000000000000000000000000000000" , -- ADDR 3641
			"00000000000000000000000000000000" , -- ADDR 3642
			"00000000000000000000000000000000" , -- ADDR 3643
			"00000000000000000000000000000000" , -- ADDR 3644
			"00000000000000000000000000000000" , -- ADDR 3645
			"00000000000000000000000000000000" , -- ADDR 3646
			"00000000000000000000000000000000" , -- ADDR 3647
			"00000000000000000000000000000000" , -- ADDR 3648
			"00000000000000000000000000000000" , -- ADDR 3649
			"00000000000000000000000000000000" , -- ADDR 3650
			"00000000000000000000000000000000" , -- ADDR 3651
			"00000000000000000000000000000000" , -- ADDR 3652
			"00000000000000000000000000000000" , -- ADDR 3653
			"00000000000000000000000000000000" , -- ADDR 3654
			"00000000000000000000000000000000" , -- ADDR 3655
			"00000000000000000000000000000000" , -- ADDR 3656
			"00000000000000000000000000000000" , -- ADDR 3657
			"00000000000000000000000000000000" , -- ADDR 3658
			"00000000000000000000000000000000" , -- ADDR 3659
			"00000000000000000000000000000000" , -- ADDR 3660
			"00000000000000000000000000000000" , -- ADDR 3661
			"00000000000000000000000000000000" , -- ADDR 3662
			"00000000000000000000000000000000" , -- ADDR 3663
			"00000000000000000000000000000000" , -- ADDR 3664
			"00000000000000000000000000000000" , -- ADDR 3665
			"00000000000000000000000000000000" , -- ADDR 3666
			"00000000000000000000000000000000" , -- ADDR 3667
			"00000000000000000000000000000000" , -- ADDR 3668
			"00000000000000000000000000000000" , -- ADDR 3669
			"00000000000000000000000000000000" , -- ADDR 3670
			"00000000000000000000000000000000" , -- ADDR 3671
			"00000000000000000000000000000000" , -- ADDR 3672
			"00000000000000000000000000000000" , -- ADDR 3673
			"00000000000000000000000000000000" , -- ADDR 3674
			"00000000000000000000000000000000" , -- ADDR 3675
			"00000000000000000000000000000000" , -- ADDR 3676
			"00000000000000000000000000000000" , -- ADDR 3677
			"00000000000000000000000000000000" , -- ADDR 3678
			"00000000000000000000000000000000" , -- ADDR 3679
			"00000000000000000000000000000000" , -- ADDR 3680
			"00000000000000000000000000000000" , -- ADDR 3681
			"00000000000000000000000000000000" , -- ADDR 3682
			"00000000000000000000000000000000" , -- ADDR 3683
			"00000000000000000000000000000000" , -- ADDR 3684
			"00000000000000000000000000000000" , -- ADDR 3685
			"00000000000000000000000000000000" , -- ADDR 3686
			"00000000000000000000000000000000" , -- ADDR 3687
			"00000000000000000000000000000000" , -- ADDR 3688
			"00000000000000000000000000000000" , -- ADDR 3689
			"00000000000000000000000000000000" , -- ADDR 3690
			"00000000000000000000000000000000" , -- ADDR 3691
			"00000000000000000000000000000000" , -- ADDR 3692
			"00000000000000000000000000000000" , -- ADDR 3693
			"00000000000000000000000000000000" , -- ADDR 3694
			"00000000000000000000000000000000" , -- ADDR 3695
			"00000000000000000000000000000000" , -- ADDR 3696
			"00000000000000000000000000000000" , -- ADDR 3697
			"00000000000000000000000000000000" , -- ADDR 3698
			"00000000000000000000000000000000" , -- ADDR 3699
			"00000000000000000000000000000000" , -- ADDR 3700
			"00000000000000000000000000000000" , -- ADDR 3701
			"00000000000000000000000000000000" , -- ADDR 3702
			"00000000000000000000000000000000" , -- ADDR 3703
			"00000000000000000000000000000000" , -- ADDR 3704
			"00000000000000000000000000000000" , -- ADDR 3705
			"00000000000000000000000000000000" , -- ADDR 3706
			"00000000000000000000000000000000" , -- ADDR 3707
			"00000000000000000000000000000000" , -- ADDR 3708
			"00000000000000000000000000000000" , -- ADDR 3709
			"00000000000000000000000000000000" , -- ADDR 3710
			"00000000000000000000000000000000" , -- ADDR 3711
			"00000000000000000000000000000000" , -- ADDR 3712
			"00000000000000000000000000000000" , -- ADDR 3713
			"00000000000000000000000000000000" , -- ADDR 3714
			"00000000000000000000000000000000" , -- ADDR 3715
			"00000000000000000000000000000000" , -- ADDR 3716
			"00000000000000000000000000000000" , -- ADDR 3717
			"00000000000000000000000000000000" , -- ADDR 3718
			"00000000000000000000000000000000" , -- ADDR 3719
			"00000000000000000000000000000000" , -- ADDR 3720
			"00000000000000000000000000000000" , -- ADDR 3721
			"00000000000000000000000000000000" , -- ADDR 3722
			"00000000000000000000000000000000" , -- ADDR 3723
			"00000000000000000000000000000000" , -- ADDR 3724
			"00000000000000000000000000000000" , -- ADDR 3725
			"00000000000000000000000000000000" , -- ADDR 3726
			"00000000000000000000000000000000" , -- ADDR 3727
			"00000000000000000000000000000000" , -- ADDR 3728
			"00000000000000000000000000000000" , -- ADDR 3729
			"00000000000000000000000000000000" , -- ADDR 3730
			"00000000000000000000000000000000" , -- ADDR 3731
			"00000000000000000000000000000000" , -- ADDR 3732
			"00000000000000000000000000000000" , -- ADDR 3733
			"00000000000000000000000000000000" , -- ADDR 3734
			"00000000000000000000000000000000" , -- ADDR 3735
			"00000000000000000000000000000000" , -- ADDR 3736
			"00000000000000000000000000000000" , -- ADDR 3737
			"00000000000000000000000000000000" , -- ADDR 3738
			"00000000000000000000000000000000" , -- ADDR 3739
			"00000000000000000000000000000000" , -- ADDR 3740
			"00000000000000000000000000000000" , -- ADDR 3741
			"00000000000000000000000000000000" , -- ADDR 3742
			"00000000000000000000000000000000" , -- ADDR 3743
			"00000000000000000000000000000000" , -- ADDR 3744
			"00000000000000000000000000000000" , -- ADDR 3745
			"00000000000000000000000000000000" , -- ADDR 3746
			"00000000000000000000000000000000" , -- ADDR 3747
			"00000000000000000000000000000000" , -- ADDR 3748
			"00000000000000000000000000000000" , -- ADDR 3749
			"00000000000000000000000000000000" , -- ADDR 3750
			"00000000000000000000000000000000" , -- ADDR 3751
			"00000000000000000000000000000000" , -- ADDR 3752
			"00000000000000000000000000000000" , -- ADDR 3753
			"00000000000000000000000000000000" , -- ADDR 3754
			"00000000000000000000000000000000" , -- ADDR 3755
			"00000000000000000000000000000000" , -- ADDR 3756
			"00000000000000000000000000000000" , -- ADDR 3757
			"00000000000000000000000000000000" , -- ADDR 3758
			"00000000000000000000000000000000" , -- ADDR 3759
			"00000000000000000000000000000000" , -- ADDR 3760
			"00000000000000000000000000000000" , -- ADDR 3761
			"00000000000000000000000000000000" , -- ADDR 3762
			"00000000000000000000000000000000" , -- ADDR 3763
			"00000000000000000000000000000000" , -- ADDR 3764
			"00000000000000000000000000000000" , -- ADDR 3765
			"00000000000000000000000000000000" , -- ADDR 3766
			"00000000000000000000000000000000" , -- ADDR 3767
			"00000000000000000000000000000000" , -- ADDR 3768
			"00000000000000000000000000000000" , -- ADDR 3769
			"00000000000000000000000000000000" , -- ADDR 3770
			"00000000000000000000000000000000" , -- ADDR 3771
			"00000000000000000000000000000000" , -- ADDR 3772
			"00000000000000000000000000000000" , -- ADDR 3773
			"00000000000000000000000000000000" , -- ADDR 3774
			"00000000000000000000000000000000" , -- ADDR 3775
			"00000000000000000000000000000000" , -- ADDR 3776
			"00000000000000000000000000000000" , -- ADDR 3777
			"00000000000000000000000000000000" , -- ADDR 3778
			"00000000000000000000000000000000" , -- ADDR 3779
			"00000000000000000000000000000000" , -- ADDR 3780
			"00000000000000000000000000000000" , -- ADDR 3781
			"00000000000000000000000000000000" , -- ADDR 3782
			"00000000000000000000000000000000" , -- ADDR 3783
			"00000000000000000000000000000000" , -- ADDR 3784
			"00000000000000000000000000000000" , -- ADDR 3785
			"00000000000000000000000000000000" , -- ADDR 3786
			"00000000000000000000000000000000" , -- ADDR 3787
			"00000000000000000000000000000000" , -- ADDR 3788
			"00000000000000000000000000000000" , -- ADDR 3789
			"00000000000000000000000000000000" , -- ADDR 3790
			"00000000000000000000000000000000" , -- ADDR 3791
			"00000000000000000000000000000000" , -- ADDR 3792
			"00000000000000000000000000000000" , -- ADDR 3793
			"00000000000000000000000000000000" , -- ADDR 3794
			"00000000000000000000000000000000" , -- ADDR 3795
			"00000000000000000000000000000000" , -- ADDR 3796
			"00000000000000000000000000000000" , -- ADDR 3797
			"00000000000000000000000000000000" , -- ADDR 3798
			"00000000000000000000000000000000" , -- ADDR 3799
			"00000000000000000000000000000000" , -- ADDR 3800
			"00000000000000000000000000000000" , -- ADDR 3801
			"00000000000000000000000000000000" , -- ADDR 3802
			"00000000000000000000000000000000" , -- ADDR 3803
			"00000000000000000000000000000000" , -- ADDR 3804
			"00000000000000000000000000000000" , -- ADDR 3805
			"00000000000000000000000000000000" , -- ADDR 3806
			"00000000000000000000000000000000" , -- ADDR 3807
			"00000000000000000000000000000000" , -- ADDR 3808
			"00000000000000000000000000000000" , -- ADDR 3809
			"00000000000000000000000000000000" , -- ADDR 3810
			"00000000000000000000000000000000" , -- ADDR 3811
			"00000000000000000000000000000000" , -- ADDR 3812
			"00000000000000000000000000000000" , -- ADDR 3813
			"00000000000000000000000000000000" , -- ADDR 3814
			"00000000000000000000000000000000" , -- ADDR 3815
			"00000000000000000000000000000000" , -- ADDR 3816
			"00000000000000000000000000000000" , -- ADDR 3817
			"00000000000000000000000000000000" , -- ADDR 3818
			"00000000000000000000000000000000" , -- ADDR 3819
			"00000000000000000000000000000000" , -- ADDR 3820
			"00000000000000000000000000000000" , -- ADDR 3821
			"00000000000000000000000000000000" , -- ADDR 3822
			"00000000000000000000000000000000" , -- ADDR 3823
			"00000000000000000000000000000000" , -- ADDR 3824
			"00000000000000000000000000000000" , -- ADDR 3825
			"00000000000000000000000000000000" , -- ADDR 3826
			"00000000000000000000000000000000" , -- ADDR 3827
			"00000000000000000000000000000000" , -- ADDR 3828
			"00000000000000000000000000000000" , -- ADDR 3829
			"00000000000000000000000000000000" , -- ADDR 3830
			"00000000000000000000000000000000" , -- ADDR 3831
			"00000000000000000000000000000000" , -- ADDR 3832
			"00000000000000000000000000000000" , -- ADDR 3833
			"00000000000000000000000000000000" , -- ADDR 3834
			"00000000000000000000000000000000" , -- ADDR 3835
			"00000000000000000000000000000000" , -- ADDR 3836
			"00000000000000000000000000000000" , -- ADDR 3837
			"00000000000000000000000000000000" , -- ADDR 3838
			"00000000000000000000000000000000" , -- ADDR 3839
			"00000000000000000000000000000000" , -- ADDR 3840
			"00000000000000000000000000000000" , -- ADDR 3841
			"00000000000000000000000000000000" , -- ADDR 3842
			"00000000000000000000000000000000" , -- ADDR 3843
			"00000000000000000000000000000000" , -- ADDR 3844
			"00000000000000000000000000000000" , -- ADDR 3845
			"00000000000000000000000000000000" , -- ADDR 3846
			"00000000000000000000000000000000" , -- ADDR 3847
			"00000000000000000000000000000000" , -- ADDR 3848
			"00000000000000000000000000000000" , -- ADDR 3849
			"00000000000000000000000000000000" , -- ADDR 3850
			"00000000000000000000000000000000" , -- ADDR 3851
			"00000000000000000000000000000000" , -- ADDR 3852
			"00000000000000000000000000000000" , -- ADDR 3853
			"00000000000000000000000000000000" , -- ADDR 3854
			"00000000000000000000000000000000" , -- ADDR 3855
			"00000000000000000000000000000000" , -- ADDR 3856
			"00000000000000000000000000000000" , -- ADDR 3857
			"00000000000000000000000000000000" , -- ADDR 3858
			"00000000000000000000000000000000" , -- ADDR 3859
			"00000000000000000000000000000000" , -- ADDR 3860
			"00000000000000000000000000000000" , -- ADDR 3861
			"00000000000000000000000000000000" , -- ADDR 3862
			"00000000000000000000000000000000" , -- ADDR 3863
			"00000000000000000000000000000000" , -- ADDR 3864
			"00000000000000000000000000000000" , -- ADDR 3865
			"00000000000000000000000000000000" , -- ADDR 3866
			"00000000000000000000000000000000" , -- ADDR 3867
			"00000000000000000000000000000000" , -- ADDR 3868
			"00000000000000000000000000000000" , -- ADDR 3869
			"00000000000000000000000000000000" , -- ADDR 3870
			"00000000000000000000000000000000" , -- ADDR 3871
			"00000000000000000000000000000000" , -- ADDR 3872
			"00000000000000000000000000000000" , -- ADDR 3873
			"00000000000000000000000000000000" , -- ADDR 3874
			"00000000000000000000000000000000" , -- ADDR 3875
			"00000000000000000000000000000000" , -- ADDR 3876
			"00000000000000000000000000000000" , -- ADDR 3877
			"00000000000000000000000000000000" , -- ADDR 3878
			"00000000000000000000000000000000" , -- ADDR 3879
			"00000000000000000000000000000000" , -- ADDR 3880
			"00000000000000000000000000000000" , -- ADDR 3881
			"00000000000000000000000000000000" , -- ADDR 3882
			"00000000000000000000000000000000" , -- ADDR 3883
			"00000000000000000000000000000000" , -- ADDR 3884
			"00000000000000000000000000000000" , -- ADDR 3885
			"00000000000000000000000000000000" , -- ADDR 3886
			"00000000000000000000000000000000" , -- ADDR 3887
			"00000000000000000000000000000000" , -- ADDR 3888
			"00000000000000000000000000000000" , -- ADDR 3889
			"00000000000000000000000000000000" , -- ADDR 3890
			"00000000000000000000000000000000" , -- ADDR 3891
			"00000000000000000000000000000000" , -- ADDR 3892
			"00000000000000000000000000000000" , -- ADDR 3893
			"00000000000000000000000000000000" , -- ADDR 3894
			"00000000000000000000000000000000" , -- ADDR 3895
			"00000000000000000000000000000000" , -- ADDR 3896
			"00000000000000000000000000000000" , -- ADDR 3897
			"00000000000000000000000000000000" , -- ADDR 3898
			"00000000000000000000000000000000" , -- ADDR 3899
			"00000000000000000000000000000000" , -- ADDR 3900
			"00000000000000000000000000000000" , -- ADDR 3901
			"00000000000000000000000000000000" , -- ADDR 3902
			"00000000000000000000000000000000" , -- ADDR 3903
			"00000000000000000000000000000000" , -- ADDR 3904
			"00000000000000000000000000000000" , -- ADDR 3905
			"00000000000000000000000000000000" , -- ADDR 3906
			"00000000000000000000000000000000" , -- ADDR 3907
			"00000000000000000000000000000000" , -- ADDR 3908
			"00000000000000000000000000000000" , -- ADDR 3909
			"00000000000000000000000000000000" , -- ADDR 3910
			"00000000000000000000000000000000" , -- ADDR 3911
			"00000000000000000000000000000000" , -- ADDR 3912
			"00000000000000000000000000000000" , -- ADDR 3913
			"00000000000000000000000000000000" , -- ADDR 3914
			"00000000000000000000000000000000" , -- ADDR 3915
			"00000000000000000000000000000000" , -- ADDR 3916
			"00000000000000000000000000000000" , -- ADDR 3917
			"00000000000000000000000000000000" , -- ADDR 3918
			"00000000000000000000000000000000" , -- ADDR 3919
			"00000000000000000000000000000000" , -- ADDR 3920
			"00000000000000000000000000000000" , -- ADDR 3921
			"00000000000000000000000000000000" , -- ADDR 3922
			"00000000000000000000000000000000" , -- ADDR 3923
			"00000000000000000000000000000000" , -- ADDR 3924
			"00000000000000000000000000000000" , -- ADDR 3925
			"00000000000000000000000000000000" , -- ADDR 3926
			"00000000000000000000000000000000" , -- ADDR 3927
			"00000000000000000000000000000000" , -- ADDR 3928
			"00000000000000000000000000000000" , -- ADDR 3929
			"00000000000000000000000000000000" , -- ADDR 3930
			"00000000000000000000000000000000" , -- ADDR 3931
			"00000000000000000000000000000000" , -- ADDR 3932
			"00000000000000000000000000000000" , -- ADDR 3933
			"00000000000000000000000000000000" , -- ADDR 3934
			"00000000000000000000000000000000" , -- ADDR 3935
			"00000000000000000000000000000000" , -- ADDR 3936
			"00000000000000000000000000000000" , -- ADDR 3937
			"00000000000000000000000000000000" , -- ADDR 3938
			"00000000000000000000000000000000" , -- ADDR 3939
			"00000000000000000000000000000000" , -- ADDR 3940
			"00000000000000000000000000000000" , -- ADDR 3941
			"00000000000000000000000000000000" , -- ADDR 3942
			"00000000000000000000000000000000" , -- ADDR 3943
			"00000000000000000000000000000000" , -- ADDR 3944
			"00000000000000000000000000000000" , -- ADDR 3945
			"00000000000000000000000000000000" , -- ADDR 3946
			"00000000000000000000000000000000" , -- ADDR 3947
			"00000000000000000000000000000000" , -- ADDR 3948
			"00000000000000000000000000000000" , -- ADDR 3949
			"00000000000000000000000000000000" , -- ADDR 3950
			"00000000000000000000000000000000" , -- ADDR 3951
			"00000000000000000000000000000000" , -- ADDR 3952
			"00000000000000000000000000000000" , -- ADDR 3953
			"00000000000000000000000000000000" , -- ADDR 3954
			"00000000000000000000000000000000" , -- ADDR 3955
			"00000000000000000000000000000000" , -- ADDR 3956
			"00000000000000000000000000000000" , -- ADDR 3957
			"00000000000000000000000000000000" , -- ADDR 3958
			"00000000000000000000000000000000" , -- ADDR 3959
			"00000000000000000000000000000000" , -- ADDR 3960
			"00000000000000000000000000000000" , -- ADDR 3961
			"00000000000000000000000000000000" , -- ADDR 3962
			"00000000000000000000000000000000" , -- ADDR 3963
			"00000000000000000000000000000000" , -- ADDR 3964
			"00000000000000000000000000000000" , -- ADDR 3965
			"00000000000000000000000000000000" , -- ADDR 3966
			"00000000000000000000000000000000" , -- ADDR 3967
			"00000000000000000000000000000000" , -- ADDR 3968
			"00000000000000000000000000000000" , -- ADDR 3969
			"00000000000000000000000000000000" , -- ADDR 3970
			"00000000000000000000000000000000" , -- ADDR 3971
			"00000000000000000000000000000000" , -- ADDR 3972
			"00000000000000000000000000000000" , -- ADDR 3973
			"00000000000000000000000000000000" , -- ADDR 3974
			"00000000000000000000000000000000" , -- ADDR 3975
			"00000000000000000000000000000000" , -- ADDR 3976
			"00000000000000000000000000000000" , -- ADDR 3977
			"00000000000000000000000000000000" , -- ADDR 3978
			"00000000000000000000000000000000" , -- ADDR 3979
			"00000000000000000000000000000000" , -- ADDR 3980
			"00000000000000000000000000000000" , -- ADDR 3981
			"00000000000000000000000000000000" , -- ADDR 3982
			"00000000000000000000000000000000" , -- ADDR 3983
			"00000000000000000000000000000000" , -- ADDR 3984
			"00000000000000000000000000000000" , -- ADDR 3985
			"00000000000000000000000000000000" , -- ADDR 3986
			"00000000000000000000000000000000" , -- ADDR 3987
			"00000000000000000000000000000000" , -- ADDR 3988
			"00000000000000000000000000000000" , -- ADDR 3989
			"00000000000000000000000000000000" , -- ADDR 3990
			"00000000000000000000000000000000" , -- ADDR 3991
			"00000000000000000000000000000000" , -- ADDR 3992
			"00000000000000000000000000000000" , -- ADDR 3993
			"00000000000000000000000000000000" , -- ADDR 3994
			"00000000000000000000000000000000" , -- ADDR 3995
			"00000000000000000000000000000000" , -- ADDR 3996
			"00000000000000000000000000000000" , -- ADDR 3997
			"00000000000000000000000000000000" , -- ADDR 3998
			"00000000000000000000000000000000" , -- ADDR 3999
			"00000000000000000000000000000000" , -- ADDR 4000
			"00000000000000000000000000000000" , -- ADDR 4001
			"00000000000000000000000000000000" , -- ADDR 4002
			"00000000000000000000000000000000" , -- ADDR 4003
			"00000000000000000000000000000000" , -- ADDR 4004
			"00000000000000000000000000000000" , -- ADDR 4005
			"00000000000000000000000000000000" , -- ADDR 4006
			"00000000000000000000000000000000" , -- ADDR 4007
			"00000000000000000000000000000000" , -- ADDR 4008
			"00000000000000000000000000000000" , -- ADDR 4009
			"00000000000000000000000000000000" , -- ADDR 4010
			"00000000000000000000000000000000" , -- ADDR 4011
			"00000000000000000000000000000000" , -- ADDR 4012
			"00000000000000000000000000000000" , -- ADDR 4013
			"00000000000000000000000000000000" , -- ADDR 4014
			"00000000000000000000000000000000" , -- ADDR 4015
			"00000000000000000000000000000000" , -- ADDR 4016
			"00000000000000000000000000000000" , -- ADDR 4017
			"00000000000000000000000000000000" , -- ADDR 4018
			"00000000000000000000000000000000" , -- ADDR 4019
			"00000000000000000000000000000000" , -- ADDR 4020
			"00000000000000000000000000000000" , -- ADDR 4021
			"00000000000000000000000000000000" , -- ADDR 4022
			"00000000000000000000000000000000" , -- ADDR 4023
			"00000000000000000000000000000000" , -- ADDR 4024
			"00000000000000000000000000000000" , -- ADDR 4025
			"00000000000000000000000000000000" , -- ADDR 4026
			"00000000000000000000000000000000" , -- ADDR 4027
			"00000000000000000000000000000000" , -- ADDR 4028
			"00000000000000000000000000000000" , -- ADDR 4029
			"00000000000000000000000000000000" , -- ADDR 4030
			"00000000000000000000000000000000" , -- ADDR 4031
			"00000000000000000000000000000000" , -- ADDR 4032
			"00000000000000000000000000000000" , -- ADDR 4033
			"00000000000000000000000000000000" , -- ADDR 4034
			"00000000000000000000000000000000" , -- ADDR 4035
			"00000000000000000000000000000000" , -- ADDR 4036
			"00000000000000000000000000000000" , -- ADDR 4037
			"00000000000000000000000000000000" , -- ADDR 4038
			"00000000000000000000000000000000" , -- ADDR 4039
			"00000000000000000000000000000000" , -- ADDR 4040
			"00000000000000000000000000000000" , -- ADDR 4041
			"00000000000000000000000000000000" , -- ADDR 4042
			"00000000000000000000000000000000" , -- ADDR 4043
			"00000000000000000000000000000000" , -- ADDR 4044
			"00000000000000000000000000000000" , -- ADDR 4045
			"00000000000000000000000000000000" , -- ADDR 4046
			"00000000000000000000000000000000" , -- ADDR 4047
			"00000000000000000000000000000000" , -- ADDR 4048
			"00000000000000000000000000000000" , -- ADDR 4049
			"00000000000000000000000000000000" , -- ADDR 4050
			"00000000000000000000000000000000" , -- ADDR 4051
			"00000000000000000000000000000000" , -- ADDR 4052
			"00000000000000000000000000000000" , -- ADDR 4053
			"00000000000000000000000000000000" , -- ADDR 4054
			"00000000000000000000000000000000" , -- ADDR 4055
			"00000000000000000000000000000000" , -- ADDR 4056
			"00000000000000000000000000000000" , -- ADDR 4057
			"00000000000000000000000000000000" , -- ADDR 4058
			"00000000000000000000000000000000" , -- ADDR 4059
			"00000000000000000000000000000000" , -- ADDR 4060
			"00000000000000000000000000000000" , -- ADDR 4061
			"00000000000000000000000000000000" , -- ADDR 4062
			"00000000000000000000000000000000" , -- ADDR 4063
			"00000000000000000000000000000000" , -- ADDR 4064
			"00000000000000000000000000000000" , -- ADDR 4065
			"00000000000000000000000000000000" , -- ADDR 4066
			"00000000000000000000000000000000" , -- ADDR 4067
			"00000000000000000000000000000000" , -- ADDR 4068
			"00000000000000000000000000000000" , -- ADDR 4069
			"00000000000000000000000000000000" , -- ADDR 4070
			"00000000000000000000000000000000" , -- ADDR 4071
			"00000000000000000000000000000000" , -- ADDR 4072
			"00000000000000000000000000000000" , -- ADDR 4073
			"00000000000000000000000000000000" , -- ADDR 4074
			"00000000000000000000000000000000" , -- ADDR 4075
			"00000000000000000000000000000000" , -- ADDR 4076
			"00000000000000000000000000000000" , -- ADDR 4077
			"00000000000000000000000000000000" , -- ADDR 4078
			"00000000000000000000000000000000" , -- ADDR 4079
			"00000000000000000000000000000000" , -- ADDR 4080
			"00000000000000000000000000000000" , -- ADDR 4081
			"00000000000000000000000000000000" , -- ADDR 4082
			"00000000000000000000000000000000" , -- ADDR 4083
			"00000000000000000000000000000000" , -- ADDR 4084
			"00000000000000000000000000000000" , -- ADDR 4085
			"00000000000000000000000000000000" , -- ADDR 4086
			"00000000000000000000000000000000" , -- ADDR 4087
			"00000000000000000000000000000000" , -- ADDR 4088
			"00000000000000000000000000000000" , -- ADDR 4089
			"00000000000000000000000000000000" , -- ADDR 4090
			"00000000000000000000000000000000" , -- ADDR 4091
			"00000000000000000000000000000000" , -- ADDR 4092
			"00000000000000000000000000000000" , -- ADDR 4093
			"00000000000000000000000000000000" , -- ADDR 4094
			"00000000000000000000000000000000"   -- ADDR 4095
			);
			
begin
	
	process (CLK)
	begin
		if (rising_edge(CLK)) then
			-- In the case of Altera Quartus, it is extremely essential that the output assignment stays in the process.
			-- Otherwise, Altera Quartus will not infer the VHDL code as ROM.
			-- However, in the case of Xilinx ISE, it does not matter whether the output assignment stays in the process
			-- or outside of it with synchronization to the clock pulse by another signal. The VHDL code will infer as ROM anyway.
			DATA <= ROM (to_integer(unsigned(ADDR)));
		end if;
	end process;
	
end Behavioral;

-- Extremely important: In order for Altera Quartus to infer the VHDL code as ROM, the setting in the path
-- "Assignments/Device…/Device and Pin Options…/Configuration/Configuration mode" must be changed to
-- "Single Uncompressed Image with memory initialization (512 Kbits UFM)".
